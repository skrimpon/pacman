module pacman_eatghost6(in, out, clk); //ok
 input [9:0] in;
 input clk;
 output reg [8:0] out;
 
 reg  [8:0] mem [0:387];
 always @(posedge clk) out  =  mem[ in ];
 
 initial begin
		mem[  0] = 9'd3;
		mem[  1] = 9'd230;
		mem[  2] = 9'd327;
		mem[  3] = 9'd245;
		mem[  4] = 9'd157;
		mem[  5] = 9'd157;
		mem[  6] = 9'd125;
		mem[  7] = 9'd117;
		mem[  8] = 9'd118;
		mem[  9] = 9'd100;
		mem[ 10] = 9'd95;
		mem[ 11] = 9'd94;
		mem[ 12] = 9'd94;
		mem[ 13] = 9'd80;
		mem[ 14] = 9'd79;
		mem[ 15] = 9'd79;
		mem[ 16] = 9'd78;
		mem[ 17] = 9'd76;
		mem[ 18] = 9'd67;
		mem[ 19] = 9'd67;
		mem[ 20] = 9'd67;
		mem[ 21] = 9'd68;
		mem[ 22] = 9'd67;
		mem[ 23] = 9'd60;
		mem[ 24] = 9'd59;
		mem[ 25] = 9'd59;
		mem[ 26] = 9'd59;
		mem[ 27] = 9'd59;
		mem[ 28] = 9'd59;
		mem[ 29] = 9'd55;
		mem[ 30] = 9'd52;
		mem[ 31] = 9'd53;
		mem[ 32] = 9'd52;
		mem[ 33] = 9'd52;
		mem[ 34] = 9'd52;
		mem[ 35] = 9'd52;
		mem[ 36] = 9'd49;
		mem[ 37] = 9'd47;
		mem[ 38] = 9'd47;
		mem[ 39] = 9'd48;
		mem[ 40] = 9'd46;
		mem[ 41] = 9'd48;
		mem[ 42] = 9'd47;
		mem[ 43] = 9'd47;
		mem[ 44] = 9'd43;
		mem[ 45] = 9'd43;
		mem[ 46] = 9'd43;
		mem[ 47] = 9'd43;
		mem[ 48] = 9'd43;
		mem[ 49] = 9'd43;
		mem[ 50] = 9'd42;
		mem[ 51] = 9'd43;
		mem[ 52] = 9'd41;
		mem[ 53] = 9'd39;
		mem[ 54] = 9'd39;
		mem[ 55] = 9'd40;
		mem[ 56] = 9'd39;
		mem[ 57] = 9'd39;
		mem[ 58] = 9'd40;
		mem[ 59] = 9'd39;
		mem[ 60] = 9'd39;
		mem[ 61] = 9'd39;
		mem[ 62] = 9'd36;
		mem[ 63] = 9'd37;
		mem[ 64] = 9'd37;
		mem[ 65] = 9'd36;
		mem[ 66] = 9'd35;
		mem[ 67] = 9'd36;
		mem[ 68] = 9'd36;
		mem[ 69] = 9'd37;
		mem[ 70] = 9'd36;
		mem[ 71] = 9'd36;
		mem[ 72] = 9'd33;
		mem[ 73] = 9'd34;
		mem[ 74] = 9'd34;
		mem[ 75] = 9'd34;
		mem[ 76] = 9'd33;
		mem[ 77] = 9'd34;
		mem[ 78] = 9'd34;
		mem[ 79] = 9'd34;
		mem[ 80] = 9'd34;
		mem[ 81] = 9'd33;
		mem[ 82] = 9'd32;
		mem[ 83] = 9'd32;
		mem[ 84] = 9'd31;
		mem[ 85] = 9'd32;
		mem[ 86] = 9'd31;
		mem[ 87] = 9'd31;
		mem[ 88] = 9'd32;
		mem[ 89] = 9'd31;
		mem[ 90] = 9'd32;
		mem[ 91] = 9'd31;
		mem[ 92] = 9'd32;
		mem[ 93] = 9'd31;
		mem[ 94] = 9'd30;
		mem[ 95] = 9'd30;
		mem[ 96] = 9'd30;
		mem[ 97] = 9'd29;
		mem[ 98] = 9'd29;
		mem[ 99] = 9'd29;
		mem[   100] = 9'd29;
		mem[   101] = 9'd30;
		mem[   102] = 9'd29;
		mem[   103] = 9'd30;
		mem[   104] = 9'd29;
		mem[   105] = 9'd30;
		mem[   106] = 9'd29;
		mem[   107] = 9'd27;
		mem[   108] = 9'd28;
		mem[   109] = 9'd28;
		mem[   110] = 9'd28;
		mem[   111] = 9'd28;
		mem[   112] = 9'd28;
		mem[   113] = 9'd27;
		mem[   114] = 9'd27;
		mem[   115] = 9'd28;
		mem[   116] = 9'd28;
		mem[   117] = 9'd27;
		mem[   118] = 9'd28;
		mem[   119] = 9'd28;
		mem[   120] = 9'd26;
		mem[   121] = 9'd26;
		mem[   122] = 9'd26;
		mem[   123] = 9'd26;
		mem[   124] = 9'd27;
		mem[   125] = 9'd26;
		mem[   126] = 9'd26;
		mem[   127] = 9'd26;
		mem[   128] = 9'd27;
		mem[   129] = 9'd26;
		mem[   130] = 9'd26;
		mem[   131] = 9'd26;
		mem[   132] = 9'd26;
		mem[   133] = 9'd26;
		mem[   134] = 9'd24;
		mem[   135] = 9'd25;
		mem[   136] = 9'd25;
		mem[   137] = 9'd25;
		mem[   138] = 9'd25;
		mem[   139] = 9'd24;
		mem[   140] = 9'd25;
		mem[   141] = 9'd25;
		mem[   142] = 9'd25;
		mem[   143] = 9'd25;
		mem[   144] = 9'd25;
		mem[   145] = 9'd25;
		mem[   146] = 9'd24;
		mem[   147] = 9'd25;
		mem[   148] = 9'd24;
		mem[   149] = 9'd23;
		mem[   150] = 9'd24;
		mem[   151] = 9'd23;
		mem[   152] = 9'd24;
		mem[   153] = 9'd24;
		mem[   154] = 9'd23;
		mem[   155] = 9'd24;
		mem[   156] = 9'd23;
		mem[   157] = 9'd24;
		mem[   158] = 9'd24;
		mem[   159] = 9'd23;
		mem[   160] = 9'd25;
		mem[   161] = 9'd23;
		mem[   162] = 9'd23;
		mem[   163] = 9'd23;
		mem[   164] = 9'd22;
		mem[   165] = 9'd23;
		mem[   166] = 9'd22;
		mem[   167] = 9'd23;
		mem[   168] = 9'd22;
		mem[   169] = 9'd22;
		mem[   170] = 9'd23;
		mem[   171] = 9'd22;
		mem[   172] = 9'd23;
		mem[   173] = 9'd23;
		mem[   174] = 9'd22;
		mem[   175] = 9'd23;
		mem[   176] = 9'd23;
		mem[   177] = 9'd22;
		mem[   178] = 9'd22;
		mem[   179] = 9'd22;
		mem[   180] = 9'd22;
		mem[   181] = 9'd21;
		mem[   182] = 9'd21;
		mem[   183] = 9'd22;
		mem[   184] = 9'd21;
		mem[   185] = 9'd21;
		mem[   186] = 9'd22;
		mem[   187] = 9'd21;
		mem[   188] = 9'd22;
		mem[   189] = 9'd21;
		mem[   190] = 9'd22;
		mem[   191] = 9'd21;
		mem[   192] = 9'd22;
		mem[   193] = 9'd22;
		mem[   194] = 9'd20;
		mem[   195] = 9'd22;
		mem[   196] = 9'd21;
		mem[   197] = 9'd21;
		mem[   198] = 9'd20;
		mem[   199] = 9'd21;
		mem[   200] = 9'd20;
		mem[   201] = 9'd20;
		mem[   202] = 9'd21;
		mem[   203] = 9'd21;
		mem[   204] = 9'd20;
		mem[   205] = 9'd21;
		mem[   206] = 9'd20;
		mem[   207] = 9'd21;
		mem[   208] = 9'd21;
		mem[   209] = 9'd20;
		mem[   210] = 9'd20;
		mem[   211] = 9'd20;
		mem[   212] = 9'd21;
		mem[   213] = 9'd20;
		mem[   214] = 9'd21;
		mem[   215] = 9'd19;
		mem[   216] = 9'd20;
		mem[   217] = 9'd20;
		mem[   218] = 9'd19;
		mem[   219] = 9'd20;
		mem[   220] = 9'd20;
		mem[   221] = 9'd19;
		mem[   222] = 9'd20;
		mem[   223] = 9'd20;
		mem[   224] = 9'd20;
		mem[   225] = 9'd19;
		mem[   226] = 9'd20;
		mem[   227] = 9'd19;
		mem[   228] = 9'd20;
		mem[   229] = 9'd19;
		mem[   230] = 9'd20;
		mem[   231] = 9'd19;
		mem[   232] = 9'd20;
		mem[   233] = 9'd19;
		mem[   234] = 9'd19;
		mem[   235] = 9'd19;
		mem[   236] = 9'd19;
		mem[   237] = 9'd19;
		mem[   238] = 9'd19;
		mem[   239] = 9'd19;
		mem[   240] = 9'd19;
		mem[   241] = 9'd19;
		mem[   242] = 9'd18;
		mem[   243] = 9'd19;
		mem[   244] = 9'd18;
		mem[   245] = 9'd19;
		mem[   246] = 9'd19;
		mem[   247] = 9'd19;
		mem[   248] = 9'd19;
		mem[   249] = 9'd19;
		mem[   250] = 9'd19;
		mem[   251] = 9'd19;
		mem[   252] = 9'd18;
		mem[   253] = 9'd18;
		mem[   254] = 9'd19;
		mem[   255] = 9'd18;
		mem[   256] = 9'd19;
		mem[   257] = 9'd17;
		mem[   258] = 9'd18;
		mem[   259] = 9'd18;
		mem[   260] = 9'd18;
		mem[   261] = 9'd18;
		mem[   262] = 9'd18;
		mem[   263] = 9'd18;
		mem[   264] = 9'd18;
		mem[   265] = 9'd18;
		mem[   266] = 9'd19;
		mem[   267] = 9'd18;
		mem[   268] = 9'd18;
		mem[   269] = 9'd19;
		mem[   270] = 9'd18;
		mem[   271] = 9'd18;
		mem[   272] = 9'd19;
		mem[   273] = 9'd17;
		mem[   274] = 9'd17;
		mem[   275] = 9'd17;
		mem[   276] = 9'd17;
		mem[   277] = 9'd18;
		mem[   278] = 9'd17;
		mem[   279] = 9'd18;
		mem[   280] = 9'd17;
		mem[   281] = 9'd17;
		mem[   282] = 9'd18;
		mem[   283] = 9'd17;
		mem[   284] = 9'd18;
		mem[   285] = 9'd17;
		mem[   286] = 9'd18;
		mem[   287] = 9'd18;
		mem[   288] = 9'd17;
		mem[   289] = 9'd18;
		mem[   290] = 9'd17;
		mem[   291] = 9'd17;
		mem[   292] = 9'd18;
		mem[   293] = 9'd17;
		mem[   294] = 9'd17;
		mem[   295] = 9'd16;
		mem[   296] = 9'd17;
		mem[   297] = 9'd17;
		mem[   298] = 9'd17;
		mem[   299] = 9'd17;
		mem[   300] = 9'd17;
		mem[   301] = 9'd17;
		mem[   302] = 9'd16;
		mem[   303] = 9'd17;
		mem[   304] = 9'd18;
		mem[   305] = 9'd16;
		mem[   306] = 9'd17;
		mem[   307] = 9'd16;
		mem[   308] = 9'd17;
		mem[   309] = 9'd17;
		mem[   310] = 9'd17;
		mem[   311] = 9'd17;
		mem[   312] = 9'd16;
		mem[   313] = 9'd17;
		mem[   314] = 9'd17;
		mem[   315] = 9'd17;
		mem[   316] = 9'd16;
		mem[   317] = 9'd16;
		mem[   318] = 9'd17;
		mem[   319] = 9'd16;
		mem[   320] = 9'd16;
		mem[   321] = 9'd17;
		mem[   322] = 9'd16;
		mem[   323] = 9'd16;
		mem[   324] = 9'd16;
		mem[   325] = 9'd16;
		mem[   326] = 9'd16;
		mem[   327] = 9'd16;
		mem[   328] = 9'd16;
		mem[   329] = 9'd17;
		mem[   330] = 9'd16;
		mem[   331] = 9'd16;
		mem[   332] = 9'd17;
		mem[   333] = 9'd16;
		mem[   334] = 9'd16;
		mem[   335] = 9'd17;
		mem[   336] = 9'd17;
		mem[   337] = 9'd16;
		mem[   338] = 9'd15;
		mem[   339] = 9'd15;
		mem[   340] = 9'd16;
		mem[   341] = 9'd16;
		mem[   342] = 9'd15;
		mem[   343] = 9'd16;
		mem[   344] = 9'd16;
		mem[   345] = 9'd15;
		mem[   346] = 9'd16;
		mem[   347] = 9'd16;
		mem[   348] = 9'd16;
		mem[   349] = 9'd15;
		mem[   350] = 9'd16;
		mem[   351] = 9'd16;
		mem[   352] = 9'd16;
		mem[   353] = 9'd15;
		mem[   354] = 9'd16;
		mem[   355] = 9'd16;
		mem[   356] = 9'd15;
		mem[   357] = 9'd16;
		mem[   358] = 9'd16;
		mem[   359] = 9'd15;
		mem[   360] = 9'd16;
		mem[   361] = 9'd15;
		mem[   362] = 9'd16;
		mem[   363] = 9'd15;
		mem[   364] = 9'd15;
		mem[   365] = 9'd15;
		mem[   366] = 9'd15;
		mem[   367] = 9'd16;
		mem[   368] = 9'd15;
		mem[   369] = 9'd15;
		mem[   370] = 9'd15;
		mem[   371] = 9'd15;
		mem[   372] = 9'd15;
		mem[   373] = 9'd16;
		mem[   374] = 9'd15;
		mem[   375] = 9'd15;
		mem[   376] = 9'd15;
		mem[   377] = 9'd15;
		mem[   378] = 9'd16;
		mem[   379] = 9'd15;
		mem[   380] = 9'd15;
		mem[   381] = 9'd15;
		mem[   382] = 9'd16;
		mem[   383] = 9'd15;
		mem[   384] = 9'd16;
		mem[   385] =  9'd511;
		mem[   386] =  9'd511;
		mem[   387] =  9'd511;
	end
	
endmodule
