module pacman_extrapac6(in, out, clk);  //ok
 input [10:0] in;
 input clk;
 output reg [8:0] out;
 
 reg  [8:0] mem [0:1096];
 always @(posedge clk) out  =  mem[ in ];
 
 initial begin
	mem[  0] = 9'd26;
	mem[  1] = 9'd44;
	mem[  2] = 9'd30;
	mem[  3] = 9'd28;
	mem[  4] = 9'd29;
	mem[  5] = 9'd29;
	mem[  6] = 9'd30;
	mem[  7] = 9'd29;
	mem[  8] = 9'd30;
	mem[  9] = 9'd29;
	mem[ 10] = 9'd29;
	mem[ 11] = 9'd30;
	mem[ 12] = 9'd59;
	mem[ 13] = 9'd58;
	mem[ 14] = 9'd30;
	mem[ 15] = 9'd29;
	mem[ 16] = 9'd30;
	mem[ 17] = 9'd29;
	mem[ 18] = 9'd30;
	mem[ 19] = 9'd29;
	mem[ 20] = 9'd30;
	mem[ 21] = 9'd29;
	mem[ 22] = 9'd29;
	mem[ 23] = 9'd30;
	mem[ 24] = 9'd29;
	mem[ 25] = 9'd30;
	mem[ 26] = 9'd29;
	mem[ 27] = 9'd30;
	mem[ 28] = 9'd29;
	mem[ 29] = 9'd30;
	mem[ 30] = 9'd29;
	mem[ 31] = 9'd30;
	mem[ 32] = 9'd29;
	mem[ 33] = 9'd29;
	mem[ 34] = 9'd30;
	mem[ 35] = 9'd29;
	mem[ 36] = 9'd30;
	mem[ 37] = 9'd29;
	mem[ 38] = 9'd30;
	mem[ 39] = 9'd29;
	mem[ 40] = 9'd30;
	mem[ 41] = 9'd29;
	mem[ 42] = 9'd30;
	mem[ 43] = 9'd29;
	mem[ 44] = 9'd29;
	mem[ 45] = 9'd30;
	mem[ 46] = 9'd29;
	mem[ 47] = 9'd30;
	mem[ 48] = 9'd29;
	mem[ 49] = 9'd30;
	mem[ 50] = 9'd29;
	mem[ 51] = 9'd29;
	mem[ 52] = 9'd30;
	mem[ 53] = 9'd29;
	mem[ 54] = 9'd30;
	mem[ 55] = 9'd29;
	mem[ 56] = 9'd30;
	mem[ 57] = 9'd29;
	mem[ 58] = 9'd30;
	mem[ 59] = 9'd29;
	mem[ 60] = 9'd29;
	mem[ 61] = 9'd30;
	mem[ 62] = 9'd29;
	mem[ 63] = 9'd30;
	mem[ 64] = 9'd29;
	mem[ 65] = 9'd30;
	mem[ 66] = 9'd29;
	mem[ 67] = 9'd30;
	mem[ 68] = 9'd29;
	mem[ 69] = 9'd29;
	mem[ 70] = 9'd30;
	mem[ 71] = 9'd29;
	mem[ 72] = 9'd30;
	mem[ 73] = 9'd29;
	mem[ 74] = 9'd30;
	mem[ 75] = 9'd29;
	mem[ 76] = 9'd30;
	mem[ 77] = 9'd29;
	mem[ 78] = 9'd30;
	mem[ 79] = 9'd29;
	mem[ 80] = 9'd29;
	mem[ 81] = 9'd30;
	mem[ 82] = 9'd29;
	mem[ 83] = 9'd30;
	mem[ 84] = 9'd58;
	mem[ 85] = 9'd59;
	mem[ 86] = 9'd59;
	mem[ 87] = 9'd59;
	mem[ 88] = 9'd59;
	mem[ 89] = 9'd59;
	mem[ 90] = 9'd59;
	mem[ 91] = 9'd59;
	mem[ 92] = 9'd58;
	mem[ 93] = 9'd59;
	mem[ 94] = 9'd59;
	mem[ 95] = 9'd59;
	mem[ 96] = 9'd59;
	mem[ 97] = 9'd59;
	mem[ 98] = 9'd59;
	mem[ 99] = 9'd59;
	mem[   100] = 9'd59;
	mem[   101] = 9'd58;
	mem[   102] = 9'd59;
	mem[   103] = 9'd59;
	mem[   104] = 9'd59;
	mem[   105] = 9'd59;
	mem[   106] = 9'd59;
	mem[   107] = 9'd59;
	mem[   108] = 9'd59;
	mem[   109] = 9'd14;
	mem[   110] = 9'd45;
	mem[   111] = 9'd29;
	mem[   112] = 9'd29;
	mem[   113] = 9'd30;
	mem[   114] = 9'd29;
	mem[   115] = 9'd29;
	mem[   116] = 9'd30;
	mem[   117] = 9'd29;
	mem[   118] = 9'd29;
	mem[   119] = 9'd30;
	mem[   120] = 9'd29;
	mem[   121] = 9'd30;
	mem[   122] = 9'd29;
	mem[   123] = 9'd30;
	mem[   124] = 9'd29;
	mem[   125] = 9'd30;
	mem[   126] = 9'd29;
	mem[   127] = 9'd30;
	mem[   128] = 9'd29;
	mem[   129] = 9'd29;
	mem[   130] = 9'd30;
	mem[   131] = 9'd29;
	mem[   132] = 9'd30;
	mem[   133] = 9'd29;
	mem[   134] = 9'd30;
	mem[   135] = 9'd29;
	mem[   136] = 9'd29;
	mem[   137] = 9'd30;
	mem[   138] = 9'd29;
	mem[   139] = 9'd30;
	mem[   140] = 9'd29;
	mem[   141] = 9'd30;
	mem[   142] = 9'd29;
	mem[   143] = 9'd30;
	mem[   144] = 9'd29;
	mem[   145] = 9'd30;
	mem[   146] = 9'd29;
	mem[   147] = 9'd30;
	mem[   148] = 9'd29;
	mem[   149] = 9'd29;
	mem[   150] = 9'd30;
	mem[   151] = 9'd29;
	mem[   152] = 9'd30;
	mem[   153] = 9'd29;
	mem[   154] = 9'd29;
	mem[   155] = 9'd30;
	mem[   156] = 9'd29;
	mem[   157] = 9'd30;
	mem[   158] = 9'd29;
	mem[   159] = 9'd30;
	mem[   160] = 9'd29;
	mem[   161] = 9'd30;
	mem[   162] = 9'd29;
	mem[   163] = 9'd30;
	mem[   164] = 9'd29;
	mem[   165] = 9'd29;
	mem[   166] = 9'd30;
	mem[   167] = 9'd29;
	mem[   168] = 9'd30;
	mem[   169] = 9'd29;
	mem[   170] = 9'd29;
	mem[   171] = 9'd30;
	mem[   172] = 9'd29;
	mem[   173] = 9'd30;
	mem[   174] = 9'd29;
	mem[   175] = 9'd30;
	mem[   176] = 9'd29;
	mem[   177] = 9'd30;
	mem[   178] = 9'd29;
	mem[   179] = 9'd30;
	mem[   180] = 9'd29;
	mem[   181] = 9'd29;
	mem[   182] = 9'd30;
	mem[   183] = 9'd59;
	mem[   184] = 9'd29;
	mem[   185] = 9'd29;
	mem[   186] = 9'd30;
	mem[   187] = 9'd29;
	mem[   188] = 9'd30;
	mem[   189] = 9'd29;
	mem[   190] = 9'd30;
	mem[   191] = 9'd29;
	mem[   192] = 9'd30;
	mem[   193] = 9'd29;
	mem[   194] = 9'd59;
	mem[   195] = 9'd59;
	mem[   196] = 9'd59;
	mem[   197] = 9'd59;
	mem[   198] = 9'd58;
	mem[   199] = 9'd59;
	mem[   200] = 9'd59;
	mem[   201] = 9'd59;
	mem[   202] = 9'd59;
	mem[   203] = 9'd59;
	mem[   204] = 9'd59;
	mem[   205] = 9'd59;
	mem[   206] = 9'd58;
	mem[   207] = 9'd59;
	mem[   208] = 9'd59;
	mem[   209] = 9'd59;
	mem[   210] = 9'd59;
	mem[   211] = 9'd59;
	mem[   212] = 9'd58;
	mem[   213] = 9'd59;
	mem[   214] = 9'd60;
	mem[   215] = 9'd58;
	mem[   216] = 9'd59;
	mem[   217] = 9'd59;
	mem[   218] = 9'd59;
	mem[   219] = 9'd385;
	mem[   220] = 9'd44;
	mem[   221] = 9'd30;
	mem[   222] = 9'd28;
	mem[   223] = 9'd29;
	mem[   224] = 9'd29;
	mem[   225] = 9'd30;
	mem[   226] = 9'd29;
	mem[   227] = 9'd30;
	mem[   228] = 9'd29;
	mem[   229] = 9'd29;
	mem[   230] = 9'd30;
	mem[   231] = 9'd59;
	mem[   232] = 9'd58;
	mem[   233] = 9'd30;
	mem[   234] = 9'd29;
	mem[   235] = 9'd30;
	mem[   236] = 9'd29;
	mem[   237] = 9'd30;
	mem[   238] = 9'd29;
	mem[   239] = 9'd30;
	mem[   240] = 9'd29;
	mem[   241] = 9'd29;
	mem[   242] = 9'd30;
	mem[   243] = 9'd29;
	mem[   244] = 9'd30;
	mem[   245] = 9'd29;
	mem[   246] = 9'd30;
	mem[   247] = 9'd29;
	mem[   248] = 9'd30;
	mem[   249] = 9'd29;
	mem[   250] = 9'd30;
	mem[   251] = 9'd29;
	mem[   252] = 9'd29;
	mem[   253] = 9'd30;
	mem[   254] = 9'd29;
	mem[   255] = 9'd30;
	mem[   256] = 9'd29;
	mem[   257] = 9'd30;
	mem[   258] = 9'd29;
	mem[   259] = 9'd30;
	mem[   260] = 9'd29;
	mem[   261] = 9'd30;
	mem[   262] = 9'd29;
	mem[   263] = 9'd29;
	mem[   264] = 9'd30;
	mem[   265] = 9'd29;
	mem[   266] = 9'd30;
	mem[   267] = 9'd29;
	mem[   268] = 9'd30;
	mem[   269] = 9'd29;
	mem[   270] = 9'd29;
	mem[   271] = 9'd30;
	mem[   272] = 9'd29;
	mem[   273] = 9'd30;
	mem[   274] = 9'd29;
	mem[   275] = 9'd30;
	mem[   276] = 9'd29;
	mem[   277] = 9'd30;
	mem[   278] = 9'd29;
	mem[   279] = 9'd29;
	mem[   280] = 9'd30;
	mem[   281] = 9'd29;
	mem[   282] = 9'd30;
	mem[   283] = 9'd29;
	mem[   284] = 9'd30;
	mem[   285] = 9'd29;
	mem[   286] = 9'd30;
	mem[   287] = 9'd29;
	mem[   288] = 9'd29;
	mem[   289] = 9'd30;
	mem[   290] = 9'd29;
	mem[   291] = 9'd30;
	mem[   292] = 9'd29;
	mem[   293] = 9'd30;
	mem[   294] = 9'd29;
	mem[   295] = 9'd30;
	mem[   296] = 9'd29;
	mem[   297] = 9'd30;
	mem[   298] = 9'd29;
	mem[   299] = 9'd29;
	mem[   300] = 9'd30;
	mem[   301] = 9'd29;
	mem[   302] = 9'd30;
	mem[   303] = 9'd58;
	mem[   304] = 9'd59;
	mem[   305] = 9'd59;
	mem[   306] = 9'd59;
	mem[   307] = 9'd59;
	mem[   308] = 9'd59;
	mem[   309] = 9'd59;
	mem[   310] = 9'd59;
	mem[   311] = 9'd58;
	mem[   312] = 9'd59;
	mem[   313] = 9'd59;
	mem[   314] = 9'd59;
	mem[   315] = 9'd59;
	mem[   316] = 9'd59;
	mem[   317] = 9'd59;
	mem[   318] = 9'd59;
	mem[   319] = 9'd59;
	mem[   320] = 9'd58;
	mem[   321] = 9'd59;
	mem[   322] = 9'd59;
	mem[   323] = 9'd59;
	mem[   324] = 9'd59;
	mem[   325] = 9'd59;
	mem[   326] = 9'd59;
	mem[   327] = 9'd59;
	mem[   328] = 9'd14;
	mem[   329] = 9'd45;
	mem[   330] = 9'd29;
	mem[   331] = 9'd29;
	mem[   332] = 9'd30;
	mem[   333] = 9'd29;
	mem[   334] = 9'd29;
	mem[   335] = 9'd30;
	mem[   336] = 9'd29;
	mem[   337] = 9'd29;
	mem[   338] = 9'd30;
	mem[   339] = 9'd29;
	mem[   340] = 9'd30;
	mem[   341] = 9'd29;
	mem[   342] = 9'd30;
	mem[   343] = 9'd29;
	mem[   344] = 9'd30;
	mem[   345] = 9'd29;
	mem[   346] = 9'd30;
	mem[   347] = 9'd29;
	mem[   348] = 9'd29;
	mem[   349] = 9'd30;
	mem[   350] = 9'd29;
	mem[   351] = 9'd30;
	mem[   352] = 9'd29;
	mem[   353] = 9'd30;
	mem[   354] = 9'd29;
	mem[   355] = 9'd29;
	mem[   356] = 9'd30;
	mem[   357] = 9'd29;
	mem[   358] = 9'd30;
	mem[   359] = 9'd29;
	mem[   360] = 9'd30;
	mem[   361] = 9'd29;
	mem[   362] = 9'd30;
	mem[   363] = 9'd29;
	mem[   364] = 9'd30;
	mem[   365] = 9'd29;
	mem[   366] = 9'd30;
	mem[   367] = 9'd29;
	mem[   368] = 9'd29;
	mem[   369] = 9'd30;
	mem[   370] = 9'd29;
	mem[   371] = 9'd30;
	mem[   372] = 9'd29;
	mem[   373] = 9'd29;
	mem[   374] = 9'd30;
	mem[   375] = 9'd29;
	mem[   376] = 9'd30;
	mem[   377] = 9'd29;
	mem[   378] = 9'd30;
	mem[   379] = 9'd29;
	mem[   380] = 9'd30;
	mem[   381] = 9'd29;
	mem[   382] = 9'd30;
	mem[   383] = 9'd29;
	mem[   384] = 9'd29;
	mem[   385] = 9'd30;
	mem[   386] = 9'd29;
	mem[   387] = 9'd30;
	mem[   388] = 9'd29;
	mem[   389] = 9'd29;
	mem[   390] = 9'd30;
	mem[   391] = 9'd29;
	mem[   392] = 9'd30;
	mem[   393] = 9'd29;
	mem[   394] = 9'd30;
	mem[   395] = 9'd29;
	mem[   396] = 9'd30;
	mem[   397] = 9'd29;
	mem[   398] = 9'd30;
	mem[   399] = 9'd29;
	mem[   400] = 9'd29;
	mem[   401] = 9'd30;
	mem[   402] = 9'd59;
	mem[   403] = 9'd29;
	mem[   404] = 9'd29;
	mem[   405] = 9'd30;
	mem[   406] = 9'd29;
	mem[   407] = 9'd30;
	mem[   408] = 9'd29;
	mem[   409] = 9'd30;
	mem[   410] = 9'd29;
	mem[   411] = 9'd30;
	mem[   412] = 9'd29;
	mem[   413] = 9'd59;
	mem[   414] = 9'd59;
	mem[   415] = 9'd59;
	mem[   416] = 9'd59;
	mem[   417] = 9'd58;
	mem[   418] = 9'd59;
	mem[   419] = 9'd59;
	mem[   420] = 9'd59;
	mem[   421] = 9'd59;
	mem[   422] = 9'd59;
	mem[   423] = 9'd59;
	mem[   424] = 9'd59;
	mem[   425] = 9'd58;
	mem[   426] = 9'd59;
	mem[   427] = 9'd59;
	mem[   428] = 9'd59;
	mem[   429] = 9'd59;
	mem[   430] = 9'd59;
	mem[   431] = 9'd58;
	mem[   432] = 9'd59;
	mem[   433] = 9'd60;
	mem[   434] = 9'd58;
	mem[   435] = 9'd59;
	mem[   436] = 9'd59;
	mem[   437] = 9'd59;
	mem[   438] = 9'd385;
	mem[   439] = 9'd44;
	mem[   440] = 9'd30;
	mem[   441] = 9'd28;
	mem[   442] = 9'd29;
	mem[   443] = 9'd29;
	mem[   444] = 9'd30;
	mem[   445] = 9'd29;
	mem[   446] = 9'd30;
	mem[   447] = 9'd29;
	mem[   448] = 9'd29;
	mem[   449] = 9'd30;
	mem[   450] = 9'd59;
	mem[   451] = 9'd58;
	mem[   452] = 9'd30;
	mem[   453] = 9'd29;
	mem[   454] = 9'd30;
	mem[   455] = 9'd29;
	mem[   456] = 9'd30;
	mem[   457] = 9'd29;
	mem[   458] = 9'd30;
	mem[   459] = 9'd29;
	mem[   460] = 9'd29;
	mem[   461] = 9'd30;
	mem[   462] = 9'd29;
	mem[   463] = 9'd30;
	mem[   464] = 9'd29;
	mem[   465] = 9'd30;
	mem[   466] = 9'd29;
	mem[   467] = 9'd30;
	mem[   468] = 9'd29;
	mem[   469] = 9'd30;
	mem[   470] = 9'd29;
	mem[   471] = 9'd29;
	mem[   472] = 9'd30;
	mem[   473] = 9'd29;
	mem[   474] = 9'd30;
	mem[   475] = 9'd29;
	mem[   476] = 9'd30;
	mem[   477] = 9'd29;
	mem[   478] = 9'd30;
	mem[   479] = 9'd29;
	mem[   480] = 9'd30;
	mem[   481] = 9'd29;
	mem[   482] = 9'd29;
	mem[   483] = 9'd30;
	mem[   484] = 9'd29;
	mem[   485] = 9'd30;
	mem[   486] = 9'd29;
	mem[   487] = 9'd30;
	mem[   488] = 9'd29;
	mem[   489] = 9'd29;
	mem[   490] = 9'd30;
	mem[   491] = 9'd29;
	mem[   492] = 9'd30;
	mem[   493] = 9'd29;
	mem[   494] = 9'd30;
	mem[   495] = 9'd29;
	mem[   496] = 9'd30;
	mem[   497] = 9'd29;
	mem[   498] = 9'd29;
	mem[   499] = 9'd30;
	mem[   500] = 9'd29;
	mem[   501] = 9'd30;
	mem[   502] = 9'd29;
	mem[   503] = 9'd30;
	mem[   504] = 9'd29;
	mem[   505] = 9'd30;
	mem[   506] = 9'd29;
	mem[   507] = 9'd29;
	mem[   508] = 9'd30;
	mem[   509] = 9'd29;
	mem[   510] = 9'd30;
	mem[   511] = 9'd29;
	mem[   512] = 9'd30;
	mem[   513] = 9'd29;
	mem[   514] = 9'd30;
	mem[   515] = 9'd29;
	mem[   516] = 9'd30;
	mem[   517] = 9'd29;
	mem[   518] = 9'd29;
	mem[   519] = 9'd30;
	mem[   520] = 9'd29;
	mem[   521] = 9'd30;
	mem[   522] = 9'd58;
	mem[   523] = 9'd59;
	mem[   524] = 9'd59;
	mem[   525] = 9'd59;
	mem[   526] = 9'd59;
	mem[   527] = 9'd59;
	mem[   528] = 9'd59;
	mem[   529] = 9'd59;
	mem[   530] = 9'd58;
	mem[   531] = 9'd59;
	mem[   532] = 9'd59;
	mem[   533] = 9'd59;
	mem[   534] = 9'd59;
	mem[   535] = 9'd59;
	mem[   536] = 9'd59;
	mem[   537] = 9'd59;
	mem[   538] = 9'd59;
	mem[   539] = 9'd58;
	mem[   540] = 9'd59;
	mem[   541] = 9'd59;
	mem[   542] = 9'd59;
	mem[   543] = 9'd59;
	mem[   544] = 9'd59;
	mem[   545] = 9'd59;
	mem[   546] = 9'd59;
	mem[   547] = 9'd14;
	mem[   548] = 9'd45;
	mem[   549] = 9'd29;
	mem[   550] = 9'd29;
	mem[   551] = 9'd30;
	mem[   552] = 9'd29;
	mem[   553] = 9'd29;
	mem[   554] = 9'd30;
	mem[   555] = 9'd29;
	mem[   556] = 9'd29;
	mem[   557] = 9'd30;
	mem[   558] = 9'd29;
	mem[   559] = 9'd30;
	mem[   560] = 9'd29;
	mem[   561] = 9'd30;
	mem[   562] = 9'd29;
	mem[   563] = 9'd30;
	mem[   564] = 9'd29;
	mem[   565] = 9'd30;
	mem[   566] = 9'd29;
	mem[   567] = 9'd29;
	mem[   568] = 9'd30;
	mem[   569] = 9'd29;
	mem[   570] = 9'd30;
	mem[   571] = 9'd29;
	mem[   572] = 9'd30;
	mem[   573] = 9'd29;
	mem[   574] = 9'd29;
	mem[   575] = 9'd30;
	mem[   576] = 9'd29;
	mem[   577] = 9'd30;
	mem[   578] = 9'd29;
	mem[   579] = 9'd30;
	mem[   580] = 9'd29;
	mem[   581] = 9'd30;
	mem[   582] = 9'd29;
	mem[   583] = 9'd30;
	mem[   584] = 9'd29;
	mem[   585] = 9'd30;
	mem[   586] = 9'd29;
	mem[   587] = 9'd29;
	mem[   588] = 9'd30;
	mem[   589] = 9'd29;
	mem[   590] = 9'd30;
	mem[   591] = 9'd29;
	mem[   592] = 9'd29;
	mem[   593] = 9'd30;
	mem[   594] = 9'd29;
	mem[   595] = 9'd30;
	mem[   596] = 9'd29;
	mem[   597] = 9'd30;
	mem[   598] = 9'd29;
	mem[   599] = 9'd30;
	mem[   600] = 9'd29;
	mem[   601] = 9'd30;
	mem[   602] = 9'd29;
	mem[   603] = 9'd29;
	mem[   604] = 9'd30;
	mem[   605] = 9'd29;
	mem[   606] = 9'd30;
	mem[   607] = 9'd29;
	mem[   608] = 9'd29;
	mem[   609] = 9'd30;
	mem[   610] = 9'd29;
	mem[   611] = 9'd30;
	mem[   612] = 9'd29;
	mem[   613] = 9'd30;
	mem[   614] = 9'd29;
	mem[   615] = 9'd30;
	mem[   616] = 9'd29;
	mem[   617] = 9'd30;
	mem[   618] = 9'd29;
	mem[   619] = 9'd29;
	mem[   620] = 9'd30;
	mem[   621] = 9'd59;
	mem[   622] = 9'd29;
	mem[   623] = 9'd29;
	mem[   624] = 9'd30;
	mem[   625] = 9'd29;
	mem[   626] = 9'd30;
	mem[   627] = 9'd29;
	mem[   628] = 9'd30;
	mem[   629] = 9'd29;
	mem[   630] = 9'd30;
	mem[   631] = 9'd29;
	mem[   632] = 9'd59;
	mem[   633] = 9'd59;
	mem[   634] = 9'd59;
	mem[   635] = 9'd59;
	mem[   636] = 9'd58;
	mem[   637] = 9'd59;
	mem[   638] = 9'd59;
	mem[   639] = 9'd59;
	mem[   640] = 9'd59;
	mem[   641] = 9'd59;
	mem[   642] = 9'd59;
	mem[   643] = 9'd59;
	mem[   644] = 9'd58;
	mem[   645] = 9'd59;
	mem[   646] = 9'd59;
	mem[   647] = 9'd59;
	mem[   648] = 9'd59;
	mem[   649] = 9'd59;
	mem[   650] = 9'd58;
	mem[   651] = 9'd59;
	mem[   652] = 9'd60;
	mem[   653] = 9'd58;
	mem[   654] = 9'd59;
	mem[   655] = 9'd59;
	mem[   656] = 9'd59;
	mem[   657] = 9'd385;
	mem[   658] = 9'd44;
	mem[   659] = 9'd30;
	mem[   660] = 9'd28;
	mem[   661] = 9'd29;
	mem[   662] = 9'd29;
	mem[   663] = 9'd30;
	mem[   664] = 9'd29;
	mem[   665] = 9'd30;
	mem[   666] = 9'd29;
	mem[   667] = 9'd29;
	mem[   668] = 9'd30;
	mem[   669] = 9'd59;
	mem[   670] = 9'd58;
	mem[   671] = 9'd30;
	mem[   672] = 9'd29;
	mem[   673] = 9'd30;
	mem[   674] = 9'd29;
	mem[   675] = 9'd30;
	mem[   676] = 9'd29;
	mem[   677] = 9'd30;
	mem[   678] = 9'd29;
	mem[   679] = 9'd29;
	mem[   680] = 9'd30;
	mem[   681] = 9'd29;
	mem[   682] = 9'd30;
	mem[   683] = 9'd29;
	mem[   684] = 9'd30;
	mem[   685] = 9'd29;
	mem[   686] = 9'd30;
	mem[   687] = 9'd29;
	mem[   688] = 9'd30;
	mem[   689] = 9'd29;
	mem[   690] = 9'd29;
	mem[   691] = 9'd30;
	mem[   692] = 9'd29;
	mem[   693] = 9'd30;
	mem[   694] = 9'd29;
	mem[   695] = 9'd30;
	mem[   696] = 9'd29;
	mem[   697] = 9'd30;
	mem[   698] = 9'd29;
	mem[   699] = 9'd30;
	mem[   700] = 9'd29;
	mem[   701] = 9'd29;
	mem[   702] = 9'd30;
	mem[   703] = 9'd29;
	mem[   704] = 9'd30;
	mem[   705] = 9'd29;
	mem[   706] = 9'd30;
	mem[   707] = 9'd29;
	mem[   708] = 9'd29;
	mem[   709] = 9'd30;
	mem[   710] = 9'd29;
	mem[   711] = 9'd30;
	mem[   712] = 9'd29;
	mem[   713] = 9'd30;
	mem[   714] = 9'd29;
	mem[   715] = 9'd30;
	mem[   716] = 9'd29;
	mem[   717] = 9'd29;
	mem[   718] = 9'd30;
	mem[   719] = 9'd29;
	mem[   720] = 9'd30;
	mem[   721] = 9'd29;
	mem[   722] = 9'd30;
	mem[   723] = 9'd29;
	mem[   724] = 9'd30;
	mem[   725] = 9'd29;
	mem[   726] = 9'd29;
	mem[   727] = 9'd30;
	mem[   728] = 9'd29;
	mem[   729] = 9'd30;
	mem[   730] = 9'd29;
	mem[   731] = 9'd30;
	mem[   732] = 9'd29;
	mem[   733] = 9'd30;
	mem[   734] = 9'd29;
	mem[   735] = 9'd30;
	mem[   736] = 9'd29;
	mem[   737] = 9'd29;
	mem[   738] = 9'd30;
	mem[   739] = 9'd29;
	mem[   740] = 9'd30;
	mem[   741] = 9'd58;
	mem[   742] = 9'd59;
	mem[   743] = 9'd59;
	mem[   744] = 9'd59;
	mem[   745] = 9'd59;
	mem[   746] = 9'd59;
	mem[   747] = 9'd59;
	mem[   748] = 9'd59;
	mem[   749] = 9'd58;
	mem[   750] = 9'd59;
	mem[   751] = 9'd59;
	mem[   752] = 9'd59;
	mem[   753] = 9'd59;
	mem[   754] = 9'd59;
	mem[   755] = 9'd59;
	mem[   756] = 9'd59;
	mem[   757] = 9'd59;
	mem[   758] = 9'd58;
	mem[   759] = 9'd59;
	mem[   760] = 9'd59;
	mem[   761] = 9'd59;
	mem[   762] = 9'd59;
	mem[   763] = 9'd59;
	mem[   764] = 9'd59;
	mem[   765] = 9'd59;
	mem[   766] = 9'd14;
	mem[   767] = 9'd45;
	mem[   768] = 9'd29;
	mem[   769] = 9'd29;
	mem[   770] = 9'd30;
	mem[   771] = 9'd29;
	mem[   772] = 9'd29;
	mem[   773] = 9'd30;
	mem[   774] = 9'd29;
	mem[   775] = 9'd29;
	mem[   776] = 9'd30;
	mem[   777] = 9'd29;
	mem[   778] = 9'd30;
	mem[   779] = 9'd29;
	mem[   780] = 9'd30;
	mem[   781] = 9'd29;
	mem[   782] = 9'd30;
	mem[   783] = 9'd29;
	mem[   784] = 9'd30;
	mem[   785] = 9'd29;
	mem[   786] = 9'd29;
	mem[   787] = 9'd30;
	mem[   788] = 9'd29;
	mem[   789] = 9'd30;
	mem[   790] = 9'd29;
	mem[   791] = 9'd30;
	mem[   792] = 9'd29;
	mem[   793] = 9'd29;
	mem[   794] = 9'd30;
	mem[   795] = 9'd29;
	mem[   796] = 9'd30;
	mem[   797] = 9'd29;
	mem[   798] = 9'd30;
	mem[   799] = 9'd29;
	mem[   800] = 9'd30;
	mem[   801] = 9'd29;
	mem[   802] = 9'd30;
	mem[   803] = 9'd29;
	mem[   804] = 9'd30;
	mem[   805] = 9'd29;
	mem[   806] = 9'd29;
	mem[   807] = 9'd30;
	mem[   808] = 9'd29;
	mem[   809] = 9'd30;
	mem[   810] = 9'd29;
	mem[   811] = 9'd29;
	mem[   812] = 9'd30;
	mem[   813] = 9'd29;
	mem[   814] = 9'd30;
	mem[   815] = 9'd29;
	mem[   816] = 9'd30;
	mem[   817] = 9'd29;
	mem[   818] = 9'd30;
	mem[   819] = 9'd29;
	mem[   820] = 9'd30;
	mem[   821] = 9'd29;
	mem[   822] = 9'd29;
	mem[   823] = 9'd30;
	mem[   824] = 9'd29;
	mem[   825] = 9'd30;
	mem[   826] = 9'd29;
	mem[   827] = 9'd29;
	mem[   828] = 9'd30;
	mem[   829] = 9'd29;
	mem[   830] = 9'd30;
	mem[   831] = 9'd29;
	mem[   832] = 9'd30;
	mem[   833] = 9'd29;
	mem[   834] = 9'd30;
	mem[   835] = 9'd29;
	mem[   836] = 9'd30;
	mem[   837] = 9'd29;
	mem[   838] = 9'd29;
	mem[   839] = 9'd30;
	mem[   840] = 9'd59;
	mem[   841] = 9'd29;
	mem[   842] = 9'd29;
	mem[   843] = 9'd30;
	mem[   844] = 9'd29;
	mem[   845] = 9'd30;
	mem[   846] = 9'd29;
	mem[   847] = 9'd30;
	mem[   848] = 9'd29;
	mem[   849] = 9'd30;
	mem[   850] = 9'd29;
	mem[   851] = 9'd59;
	mem[   852] = 9'd59;
	mem[   853] = 9'd59;
	mem[   854] = 9'd59;
	mem[   855] = 9'd58;
	mem[   856] = 9'd59;
	mem[   857] = 9'd59;
	mem[   858] = 9'd59;
	mem[   859] = 9'd59;
	mem[   860] = 9'd59;
	mem[   861] = 9'd59;
	mem[   862] = 9'd59;
	mem[   863] = 9'd58;
	mem[   864] = 9'd59;
	mem[   865] = 9'd59;
	mem[   866] = 9'd59;
	mem[   867] = 9'd59;
	mem[   868] = 9'd59;
	mem[   869] = 9'd58;
	mem[   870] = 9'd59;
	mem[   871] = 9'd60;
	mem[   872] = 9'd58;
	mem[   873] = 9'd59;
	mem[   874] = 9'd59;
	mem[   875] = 9'd59;
	mem[   876] = 9'd385;
	mem[   877] = 9'd44;
	mem[   878] = 9'd30;
	mem[   879] = 9'd28;
	mem[   880] = 9'd29;
	mem[   881] = 9'd29;
	mem[   882] = 9'd30;
	mem[   883] = 9'd29;
	mem[   884] = 9'd30;
	mem[   885] = 9'd29;
	mem[   886] = 9'd29;
	mem[   887] = 9'd30;
	mem[   888] = 9'd59;
	mem[   889] = 9'd58;
	mem[   890] = 9'd30;
	mem[   891] = 9'd29;
	mem[   892] = 9'd30;
	mem[   893] = 9'd29;
	mem[   894] = 9'd30;
	mem[   895] = 9'd29;
	mem[   896] = 9'd30;
	mem[   897] = 9'd29;
	mem[   898] = 9'd29;
	mem[   899] = 9'd30;
	mem[   900] = 9'd29;
	mem[   901] = 9'd30;
	mem[   902] = 9'd29;
	mem[   903] = 9'd30;
	mem[   904] = 9'd29;
	mem[   905] = 9'd30;
	mem[   906] = 9'd29;
	mem[   907] = 9'd30;
	mem[   908] = 9'd29;
	mem[   909] = 9'd29;
	mem[   910] = 9'd30;
	mem[   911] = 9'd29;
	mem[   912] = 9'd30;
	mem[   913] = 9'd29;
	mem[   914] = 9'd30;
	mem[   915] = 9'd29;
	mem[   916] = 9'd30;
	mem[   917] = 9'd29;
	mem[   918] = 9'd30;
	mem[   919] = 9'd29;
	mem[   920] = 9'd29;
	mem[   921] = 9'd30;
	mem[   922] = 9'd29;
	mem[   923] = 9'd30;
	mem[   924] = 9'd29;
	mem[   925] = 9'd30;
	mem[   926] = 9'd29;
	mem[   927] = 9'd29;
	mem[   928] = 9'd30;
	mem[   929] = 9'd29;
	mem[   930] = 9'd30;
	mem[   931] = 9'd29;
	mem[   932] = 9'd30;
	mem[   933] = 9'd29;
	mem[   934] = 9'd30;
	mem[   935] = 9'd29;
	mem[   936] = 9'd29;
	mem[   937] = 9'd30;
	mem[   938] = 9'd29;
	mem[   939] = 9'd30;
	mem[   940] = 9'd29;
	mem[   941] = 9'd30;
	mem[   942] = 9'd29;
	mem[   943] = 9'd30;
	mem[   944] = 9'd29;
	mem[   945] = 9'd29;
	mem[   946] = 9'd30;
	mem[   947] = 9'd29;
	mem[   948] = 9'd30;
	mem[   949] = 9'd29;
	mem[   950] = 9'd30;
	mem[   951] = 9'd29;
	mem[   952] = 9'd30;
	mem[   953] = 9'd29;
	mem[   954] = 9'd30;
	mem[   955] = 9'd29;
	mem[   956] = 9'd29;
	mem[   957] = 9'd30;
	mem[   958] = 9'd29;
	mem[   959] = 9'd30;
	mem[   960] = 9'd58;
	mem[   961] = 9'd59;
	mem[   962] = 9'd59;
	mem[   963] = 9'd59;
	mem[   964] = 9'd59;
	mem[   965] = 9'd59;
	mem[   966] = 9'd59;
	mem[   967] = 9'd59;
	mem[   968] = 9'd58;
	mem[   969] = 9'd59;
	mem[   970] = 9'd59;
	mem[   971] = 9'd59;
	mem[   972] = 9'd59;
	mem[   973] = 9'd59;
	mem[   974] = 9'd59;
	mem[   975] = 9'd59;
	mem[   976] = 9'd59;
	mem[   977] = 9'd58;
	mem[   978] = 9'd59;
	mem[   979] = 9'd59;
	mem[   980] = 9'd59;
	mem[   981] = 9'd59;
	mem[   982] = 9'd59;
	mem[   983] = 9'd59;
	mem[   984] = 9'd59;
	mem[   985] = 9'd14;
	mem[   986] = 9'd45;
	mem[   987] = 9'd29;
	mem[   988] = 9'd29;
	mem[   989] = 9'd30;
	mem[   990] = 9'd29;
	mem[   991] = 9'd29;
	mem[   992] = 9'd30;
	mem[   993] = 9'd29;
	mem[   994] = 9'd29;
	mem[   995] = 9'd30;
	mem[   996] = 9'd29;
	mem[   997] = 9'd30;
	mem[   998] = 9'd29;
	mem[   999] = 9'd30;
	mem[  1000] = 9'd29;
	mem[  1001] = 9'd30;
	mem[  1002] = 9'd29;
	mem[  1003] = 9'd30;
	mem[  1004] = 9'd29;
	mem[  1005] = 9'd29;
	mem[  1006] = 9'd30;
	mem[  1007] = 9'd29;
	mem[  1008] = 9'd30;
	mem[  1009] = 9'd29;
	mem[  1010] = 9'd30;
	mem[  1011] = 9'd29;
	mem[  1012] = 9'd29;
	mem[  1013] = 9'd30;
	mem[  1014] = 9'd29;
	mem[  1015] = 9'd30;
	mem[  1016] = 9'd29;
	mem[  1017] = 9'd30;
	mem[  1018] = 9'd29;
	mem[  1019] = 9'd30;
	mem[  1020] = 9'd29;
	mem[  1021] = 9'd30;
	mem[  1022] = 9'd29;
	mem[  1023] = 9'd30;
	mem[  1024] = 9'd29;
	mem[  1025] = 9'd29;
	mem[  1026] = 9'd30;
	mem[  1027] = 9'd29;
	mem[  1028] = 9'd30;
	mem[  1029] = 9'd29;
	mem[  1030] = 9'd29;
	mem[  1031] = 9'd30;
	mem[  1032] = 9'd29;
	mem[  1033] = 9'd30;
	mem[  1034] = 9'd29;
	mem[  1035] = 9'd30;
	mem[  1036] = 9'd29;
	mem[  1037] = 9'd30;
	mem[  1038] = 9'd29;
	mem[  1039] = 9'd30;
	mem[  1040] = 9'd29;
	mem[  1041] = 9'd29;
	mem[  1042] = 9'd30;
	mem[  1043] = 9'd29;
	mem[  1044] = 9'd30;
	mem[  1045] = 9'd29;
	mem[  1046] = 9'd29;
	mem[  1047] = 9'd30;
	mem[  1048] = 9'd29;
	mem[  1049] = 9'd30;
	mem[  1050] = 9'd29;
	mem[  1051] = 9'd30;
	mem[  1052] = 9'd29;
	mem[  1053] = 9'd30;
	mem[  1054] = 9'd29;
	mem[  1055] = 9'd30;
	mem[  1056] = 9'd29;
	mem[  1057] = 9'd29;
	mem[  1058] = 9'd30;
	mem[  1059] = 9'd59;
	mem[  1060] = 9'd29;
	mem[  1061] = 9'd29;
	mem[  1062] = 9'd30;
	mem[  1063] = 9'd29;
	mem[  1064] = 9'd30;
	mem[  1065] = 9'd29;
	mem[  1066] = 9'd30;
	mem[  1067] = 9'd29;
	mem[  1068] = 9'd30;
	mem[  1069] = 9'd29;
	mem[  1070] = 9'd59;
	mem[  1071] = 9'd59;
	mem[  1072] = 9'd59;
	mem[  1073] = 9'd59;
	mem[  1074] = 9'd58;
	mem[  1075] = 9'd59;
	mem[  1076] = 9'd59;
	mem[  1077] = 9'd59;
	mem[  1078] = 9'd59;
	mem[  1079] = 9'd59;
	mem[  1080] = 9'd59;
	mem[  1081] = 9'd59;
	mem[  1082] = 9'd58;
	mem[  1083] = 9'd59;
	mem[  1084] = 9'd59;
	mem[  1085] = 9'd59;
	mem[  1086] = 9'd59;
	mem[  1087] = 9'd59;
	mem[  1088] = 9'd58;
	mem[  1089] = 9'd59;
	mem[  1090] = 9'd60;
	mem[  1091] = 9'd58;
	mem[  1092] = 9'd59;
	mem[  1093] = 9'd59;
	mem[  1094] = 9'd59;
	mem[  1095] = 9'd511;
	mem[  1096] = 9'd511;
	end
	
endmodule

