module pacman_eatfruit6(in, out, clk); //ok
 input [6:0] in;
 input clk;
 output reg [8:0] out;
 
 reg  [8:0] mem [0:122];
 always @(posedge clk) out  =  mem[ in ];
 
 initial begin
	mem[  0] = 9'd71;
	mem[  1] = 9'd42;
	mem[  2] = 9'd41;
	mem[  3] = 9'd42;
	mem[  4] = 9'd42;
	mem[  5] = 9'd43;
	mem[  6] = 9'd42;
	mem[  7] = 9'd43;
	mem[  8] = 9'd44;
	mem[  9] = 9'd47;
	mem[ 10] = 9'd47;
	mem[ 11] = 9'd47;
	mem[ 12] = 9'd48;
	mem[ 13] = 9'd47;
	mem[ 14] = 9'd47;
	mem[ 15] = 9'd47;
	mem[ 16] = 9'd50;
	mem[ 17] = 9'd53;
	mem[ 18] = 9'd52;
	mem[ 19] = 9'd53;
	mem[ 20] = 9'd52;
	mem[ 21] = 9'd52;
	mem[ 22] = 9'd53;
	mem[ 23] = 9'd57;
	mem[ 24] = 9'd58;
	mem[ 25] = 9'd59;
	mem[ 26] = 9'd59;
	mem[ 27] = 9'd59;
	mem[ 28] = 9'd59;
	mem[ 29] = 9'd62;
	mem[ 30] = 9'd68;
	mem[ 31] = 9'd67;
	mem[ 32] = 9'd68;
	mem[ 33] = 9'd67;
	mem[ 34] = 9'd68;
	mem[ 35] = 9'd78;
	mem[ 36] = 9'd78;
	mem[ 37] = 9'd79;
	mem[ 38] = 9'd79;
	mem[ 39] = 9'd84;
	mem[ 40] = 9'd94;
	mem[ 41] = 9'd95;
	mem[ 42] = 9'd94;
	mem[ 43] = 9'd105;
	mem[ 44] = 9'd118;
	mem[ 45] = 9'd118;
	mem[ 46] = 9'd132;
	mem[ 47] = 9'd159;
	mem[ 48] = 9'd162;
	mem[ 49] = 9'd234;
	mem[ 50] = 9'd327;
	mem[ 51] = 9'd326;
	mem[ 52] = 9'd220;
	mem[ 53] = 9'd157;
	mem[ 54] = 9'd158;
	mem[ 55] = 9'd122;
	mem[ 56] = 9'd118;
	mem[ 57] = 9'd118;
	mem[ 58] = 9'd99;
	mem[ 59] = 9'd94;
	mem[ 60] = 9'd94;
	mem[ 61] = 9'd94;
	mem[ 62] = 9'd79;
	mem[ 63] = 9'd79;
	mem[ 64] = 9'd78;
	mem[ 65] = 9'd79;
	mem[ 66] = 9'd75;
	mem[ 67] = 9'd67;
	mem[ 68] = 9'd67;
	mem[ 69] = 9'd68;
	mem[ 70] = 9'd67;
	mem[ 71] = 9'd67;
	mem[ 72] = 9'd60;
	mem[ 73] = 9'd59;
	mem[ 74] = 9'd58;
	mem[ 75] = 9'd59;
	mem[ 76] = 9'd59;
	mem[ 77] = 9'd59;
	mem[ 78] = 9'd54;
	mem[ 79] = 9'd53;
	mem[ 80] = 9'd52;
	mem[ 81] = 9'd52;
	mem[ 82] = 9'd53;
	mem[ 83] = 9'd52;
	mem[ 84] = 9'd52;
	mem[ 85] = 9'd49;
	mem[ 86] = 9'd47;
	mem[ 87] = 9'd47;
	mem[ 88] = 9'd47;
	mem[ 89] = 9'd47;
	mem[ 90] = 9'd47;
	mem[ 91] = 9'd47;
	mem[ 92] = 9'd47;
	mem[ 93] = 9'd43;
	mem[ 94] = 9'd43;
	mem[ 95] = 9'd43;
	mem[ 96] = 9'd42;
	mem[ 97] = 9'd43;
	mem[ 98] = 9'd43;
	mem[ 99] = 9'd43;
	mem[   100] = 9'd43;
	mem[   101] = 9'd41;
	mem[   102] = 9'd39;
	mem[   103] = 9'd39;
	mem[   104] = 9'd39;
	mem[   105] = 9'd39;
	mem[   106] = 9'd40;
	mem[   107] = 9'd39;
	mem[   108] = 9'd39;
	mem[   109] = 9'd39;
	mem[   110] = 9'd39;
	mem[   111] = 9'd36;
	mem[   112] = 9'd36;
	mem[   113] = 9'd37;
	mem[   114] = 9'd36;
	mem[   115] = 9'd36;
	mem[   116] = 9'd36;
	mem[   117] = 9'd37;
	mem[   118] = 9'd36;
	mem[   119] = 9'd36;
	mem[   120] = 9'd30;
	mem[   121] = 9'd511;
	mem[   122] = 9'd511;
	end
	
endmodule

