module pacman_beginning_converted(in, out, clk); 
	 input [11:0] in;
	 input clk;
	 output reg [9:0] out;
	 
	 reg  [9:0] mem [0:2153];
	 always @(posedge clk) out  =  mem[ in ];
	 
	 initial begin
		mem[     0] = 10'd190;    
		mem[     1] = 10'd43;    
		mem[     2] = 10'd39;    
		mem[     3] = 10'd49;    
		mem[     4] = 10'd40;    
		mem[     5] = 10'd32;    
		mem[     6] = 10'd91;    
		mem[     7] = 10'd31;    
		mem[     8] = 10'd43;    
		mem[     9] = 10'd89;    
		mem[    10] = 10'd41;    
		mem[    11] = 10'd33;    
		mem[    12] = 10'd43;    
		mem[    13] = 10'd48;    
		mem[    14] = 10'd31;    
		mem[    15] = 10'd43;    
		mem[    16] = 10'd40;    
		mem[    17] = 10'd49;    
		mem[    18] = 10'd41;    
		mem[    19] = 10'd33;    
		mem[    20] = 10'd44;    
		mem[    21] = 10'd47;    
		mem[    22] = 10'd31;    
		mem[    23] = 10'd44;    
		mem[    24] = 10'd40;    
		mem[    25] = 10'd48;    
		mem[    26] = 10'd41;    
		mem[    27] = 10'd34;    
		mem[    28] = 10'd43;    
		mem[    29] = 10'd46;    
		mem[    30] = 10'd32;    
		mem[    31] = 10'd44;    
		mem[    32] = 10'd159;    
		mem[    33] = 10'd113;    
		mem[    34] = 10'd42;    
		mem[    35] = 10'd156;    
		mem[    36] = 10'd130;    
		mem[    37] = 10'd42;    
		mem[    38] = 10'd162;    
		mem[    39] = 10'd124;    
		mem[    40] = 10'd42;    
		mem[    41] = 10'd162;    
		mem[    42] = 10'd124;    
		mem[    43] = 10'd42;    
		mem[    44] = 10'd162;    
		mem[    45] = 10'd76;    
		mem[    46] = 10'd22;    
		mem[    47] = 10'd20;    
		mem[    48] = 10'd18;    
		mem[    49] = 10'd24;    
		mem[    50] = 10'd19;    
		mem[    51] = 10'd20;    
		mem[    52] = 10'd21;    
		mem[    53] = 10'd21;    
		mem[    54] = 10'd22;    
		mem[    55] = 10'd21;    
		mem[    56] = 10'd20;    
		mem[    57] = 10'd20;    
		mem[    58] = 10'd19;    
		mem[    59] = 10'd20;    
		mem[    60] = 10'd22;    
		mem[    61] = 10'd22;    
		mem[    62] = 10'd20;    
		mem[    63] = 10'd20;    
		mem[    64] = 10'd19;    
		mem[    65] = 10'd23;    
		mem[    66] = 10'd19;    
		mem[    67] = 10'd20;    
		mem[    68] = 10'd20;    
		mem[    69] = 10'd21;    
		mem[    70] = 10'd22;    
		mem[    71] = 10'd20;    
		mem[    72] = 10'd21;    
		mem[    73] = 10'd19;    
		mem[    74] = 10'd20;    
		mem[    75] = 10'd20;    
		mem[    76] = 10'd21;    
		mem[    77] = 10'd22;    
		mem[    78] = 10'd21;    
		mem[    79] = 10'd19;    
		mem[    80] = 10'd19;    
		mem[    81] = 10'd23;    
		mem[    82] = 10'd19;    
		mem[    83] = 10'd20;    
		mem[    84] = 10'd21;    
		mem[    85] = 10'd21;    
		mem[    86] = 10'd21;    
		mem[    87] = 10'd21;    
		mem[    88] = 10'd20;    
		mem[    89] = 10'd20;    
		mem[    90] = 10'd20;    
		mem[    91] = 10'd20;    
		mem[    92] = 10'd21;    
		mem[    93] = 10'd21;    
		mem[    94] = 10'd21;    
		mem[    95] = 10'd20;    
		mem[    96] = 10'd19;    
		mem[    97] = 10'd22;    
		mem[    98] = 10'd20;    
		mem[    99] = 10'd20;    
		mem[   100] = 10'd21;    
		mem[   101] = 10'd20;    
		mem[   102] = 10'd21;    
		mem[   103] = 10'd21;    
		mem[   104] = 10'd20;    
		mem[   105] = 10'd21;    
		mem[   106] = 10'd19;    
		mem[   107] = 10'd21;    
		mem[   108] = 10'd21;    
		mem[   109] = 10'd21;    
		mem[   110] = 10'd20;    
		mem[   111] = 10'd21;    
		mem[   112] = 10'd19;    
		mem[   113] = 10'd22;    
		mem[   114] = 10'd177;    
		mem[   115] = 10'd1023;//10'd1301;    
		mem[   116] = 10'd27;    
		mem[   117] = 10'd27;    
		mem[   118] = 10'd27;    
		mem[   119] = 10'd27;    
		mem[   120] = 10'd28;    
		mem[   121] = 10'd27;    
		mem[   122] = 10'd27;    
		mem[   123] = 10'd27;    
		mem[   124] = 10'd28;    
		mem[   125] = 10'd27;    
		mem[   126] = 10'd27;    
		mem[   127] = 10'd28;    
		mem[   128] = 10'd27;    
		mem[   129] = 10'd27;    
		mem[   130] = 10'd27;    
		mem[   131] = 10'd28;    
		mem[   132] = 10'd27;    
		mem[   133] = 10'd27;    
		mem[   134] = 10'd28;    
		mem[   135] = 10'd27;    
		mem[   136] = 10'd27;    
		mem[   137] = 10'd27;    
		mem[   138] = 10'd28;    
		mem[   139] = 10'd27;    
		mem[   140] = 10'd28;    
		mem[   141] = 10'd27;    
		mem[   142] = 10'd27;    
		mem[   143] = 10'd27;    
		mem[   144] = 10'd28;    
		mem[   145] = 10'd27;    
		mem[   146] = 10'd27;    
		mem[   147] = 10'd28;    
		mem[   148] = 10'd27;    
		mem[   149] = 10'd27;    
		mem[   150] = 10'd28;    
		mem[   151] = 10'd27;    
		mem[   152] = 10'd27;    
		mem[   153] = 10'd28;    
		mem[   154] = 10'd27;    
		mem[   155] = 10'd27;    
		mem[   156] = 10'd27;    
		mem[   157] = 10'd28;    
		mem[   158] = 10'd27;    
		mem[   159] = 10'd27;    
		mem[   160] = 10'd28;    
		mem[   161] = 10'd27;    
		mem[   162] = 10'd27;    
		mem[   163] = 10'd28;    
		mem[   164] = 10'd27;    
		mem[   165] = 10'd27;    
		mem[   166] = 10'd27;    
		mem[   167] = 10'd28;    
		mem[   168] = 10'd27;    
		mem[   169] = 10'd1023;//10'd1101;    
		mem[   170] = 10'd387;    
		mem[   171] = 10'd66;    
		mem[   172] = 10'd31;    
		mem[   173] = 10'd30;    
		mem[   174] = 10'd41;    
		mem[   175] = 10'd28;    
		mem[   176] = 10'd68;    
		mem[   177] = 10'd23;    
		mem[   178] = 10'd34;    
		mem[   179] = 10'd34;    
		mem[   180] = 10'd39;    
		mem[   181] = 10'd27;    
		mem[   182] = 10'd31;    
		mem[   183] = 10'd38;    
		mem[   184] = 10'd33;    
		mem[   185] = 10'd24;    
		mem[   186] = 10'd38;    
		mem[   187] = 10'd35;    
		mem[   188] = 10'd26;    
		mem[   189] = 10'd39;    
		mem[   190] = 10'd31;    
		mem[   191] = 10'd31;    
		mem[   192] = 10'd27;    
		mem[   193] = 10'd41;    
		mem[   194] = 10'd31;    
		mem[   195] = 10'd26;    
		mem[   196] = 10'd41;    
		mem[   197] = 10'd28;    
		mem[   198] = 10'd31;    
		mem[   199] = 10'd32;    
		mem[   200] = 10'd40;    
		mem[   201] = 10'd28;    
		mem[   202] = 10'd29;    
		mem[   203] = 10'd39;    
		mem[   204] = 10'd24;    
		mem[   205] = 10'd35;    
		mem[   206] = 10'd35;    
		mem[   207] = 10'd36;    
		mem[   208] = 10'd27;    
		mem[   209] = 10'd34;    
		mem[   210] = 10'd35;    
		mem[   211] = 10'd33;    
		mem[   212] = 10'd27;    
		mem[   213] = 10'd70;    
		mem[   214] = 10'd95;    
		mem[   215] = 10'd28;    
		mem[   216] = 10'd110;    
		mem[   217] = 10'd85;    
		mem[   218] = 10'd28;    
		mem[   219] = 10'd109;    
		mem[   220] = 10'd81;    
		mem[   221] = 10'd28;    
		mem[   222] = 10'd105;    
		mem[   223] = 10'd82;    
		mem[   224] = 10'd28;    
		mem[   225] = 10'd109;    
		mem[   226] = 10'd81;    
		mem[   227] = 10'd28;    
		mem[   228] = 10'd108;    
		mem[   229] = 10'd83;    
		mem[   230] = 10'd30;    
		mem[   231] = 10'd106;    
		mem[   232] = 10'd93;    
		mem[   233] = 10'd20;    
		mem[   234] = 10'd19;    
		mem[   235] = 10'd18;    
		mem[   236] = 10'd19;    
		mem[   237] = 10'd22;    
		mem[   238] = 10'd23;    
		mem[   239] = 10'd23;    
		mem[   240] = 10'd20;    
		mem[   241] = 10'd18;    
		mem[   242] = 10'd18;    
		mem[   243] = 10'd18;    
		mem[   244] = 10'd44;    
		mem[   245] = 10'd23;    
		mem[   246] = 10'd20;    
		mem[   247] = 10'd18;    
		mem[   248] = 10'd20;    
		mem[   249] = 10'd21;    
		mem[   250] = 10'd18;    
		mem[   251] = 10'd42;    
		mem[   252] = 10'd23;    
		mem[   253] = 10'd22;    
		mem[   254] = 10'd21;    
		mem[   255] = 10'd19;    
		mem[   256] = 10'd19;    
		mem[   257] = 10'd17;    
		mem[   258] = 10'd45;    
		mem[   259] = 10'd23;    
		mem[   260] = 10'd20;    
		mem[   261] = 10'd17;    
		mem[   262] = 10'd21;    
		mem[   263] = 10'd20;    
		mem[   264] = 10'd19;    
		mem[   265] = 10'd20;    
		mem[   266] = 10'd22;    
		mem[   267] = 10'd22;    
		mem[   268] = 10'd23;    
		mem[   269] = 10'd21;    
		mem[   270] = 10'd18;    
		mem[   271] = 10'd19;    
		mem[   272] = 10'd18;    
		mem[   273] = 10'd45;    
		mem[   274] = 10'd22;    
		mem[   275] = 10'd20;    
		mem[   276] = 10'd18;    
		mem[   277] = 10'd21;    
		mem[   278] = 10'd20;    
		mem[   279] = 10'd19;    
		mem[   280] = 10'd19;    
		mem[   281] = 10'd23;    
		mem[   282] = 10'd22;    
		mem[   283] = 10'd22;    
		mem[   284] = 10'd21;    
		mem[   285] = 10'd19;    
		mem[   286] = 10'd19;    
		mem[   287] = 10'd18;    
		mem[   288] = 10'd21;    
		mem[   289] = 10'd23;    
		mem[   290] = 10'd23;    
		mem[   291] = 10'd20;    
		mem[   292] = 10'd18;    
		mem[   293] = 10'd20;    
		mem[   294] = 10'd21;    
		mem[   295] = 10'd19;    
		mem[   296] = 10'd20;    
		mem[   297] = 10'd21;    
		mem[   298] = 10'd23;    
		mem[   299] = 10'd27;    
		mem[   300] = 10'd27;    
		mem[   301] = 10'd24;    
		mem[   302] = 10'd25;    
		mem[   303] = 10'd29;    
		mem[   304] = 10'd32;    
		mem[   305] = 10'd26;    
		mem[   306] = 10'd22;    
		mem[   307] = 10'd31;    
		mem[   308] = 10'd25;    
		mem[   309] = 10'd27;    
		mem[   310] = 10'd30;    
		mem[   311] = 10'd30;    
		mem[   312] = 10'd26;    
		mem[   313] = 10'd25;    
		mem[   314] = 10'd25;    
		mem[   315] = 10'd29;    
		mem[   316] = 10'd31;    
		mem[   317] = 10'd26;    
		mem[   318] = 10'd23;    
		mem[   319] = 10'd30;    
		mem[   320] = 10'd25;    
		mem[   321] = 10'd28;    
		mem[   322] = 10'd30;    
		mem[   323] = 10'd29;    
		mem[   324] = 10'd27;    
		mem[   325] = 10'd25;    
		mem[   326] = 10'd25;    
		mem[   327] = 10'd29;    
		mem[   328] = 10'd30;    
		mem[   329] = 10'd27;    
		mem[   330] = 10'd23;    
		mem[   331] = 10'd30;    
		mem[   332] = 10'd25;    
		mem[   333] = 10'd28;    
		mem[   334] = 10'd30;    
		mem[   335] = 10'd29;    
		mem[   336] = 10'd26;    
		mem[   337] = 10'd25;    
		mem[   338] = 10'd25;    
		mem[   339] = 10'd30;    
		mem[   340] = 10'd29;    
		mem[   341] = 10'd27;    
		mem[   342] = 10'd24;    
		mem[   343] = 10'd30;    
		mem[   344] = 10'd25;    
		mem[   345] = 10'd28;    
		mem[   346] = 10'd29;    
		mem[   347] = 10'd29;    
		mem[   348] = 10'd27;    
		mem[   349] = 10'd25;    
		mem[   350] = 10'd26;    
		mem[   351] = 10'd28;    
		mem[   352] = 10'd81;    
		mem[   353] = 10'd48;    
		mem[   354] = 10'd140;    
		mem[   355] = 10'd118;    
		mem[   356] = 10'd50;    
		mem[   357] = 10'd154;    
		mem[   358] = 10'd132;    
		mem[   359] = 10'd42;    
		mem[   360] = 10'd162;    
		mem[   361] = 10'd124;    
		mem[   362] = 10'd42;    
		mem[   363] = 10'd162;    
		mem[   364] = 10'd124;    
		mem[   365] = 10'd42;    
		mem[   366] = 10'd163;    
		mem[   367] = 10'd123;    
		mem[   368] = 10'd42;    
		mem[   369] = 10'd1023;//10'd1256;    
		mem[   370] = 10'd34;    
		mem[   371] = 10'd34;    
		mem[   372] = 10'd33;    
		mem[   373] = 10'd33;    
		mem[   374] = 10'd33;    
		mem[   375] = 10'd33;    
		mem[   376] = 10'd32;    
		mem[   377] = 10'd33;    
		mem[   378] = 10'd32;    
		mem[   379] = 10'd33;    
		mem[   380] = 10'd32;    
		mem[   381] = 10'd33;    
		mem[   382] = 10'd32;    
		mem[   383] = 10'd33;    
		mem[   384] = 10'd32;    
		mem[   385] = 10'd32;    
		mem[   386] = 10'd33;    
		mem[   387] = 10'd32;    
		mem[   388] = 10'd33;    
		mem[   389] = 10'd32;    
		mem[   390] = 10'd33;    
		mem[   391] = 10'd32;    
		mem[   392] = 10'd32;    
		mem[   393] = 10'd33;    
		mem[   394] = 10'd32;    
		mem[   395] = 10'd33;    
		mem[   396] = 10'd32;    
		mem[   397] = 10'd33;    
		mem[   398] = 10'd32;    
		mem[   399] = 10'd33;    
		mem[   400] = 10'd32;    
		mem[   401] = 10'd33;    
		mem[   402] = 10'd32;    
		mem[   403] = 10'd33;    
		mem[   404] = 10'd32;    
		mem[   405] = 10'd32;    
		mem[   406] = 10'd33;    
		mem[   407] = 10'd32;    
		mem[   408] = 10'd33;    
		mem[   409] = 10'd32;    
		mem[   410] = 10'd33;    
		mem[   411] = 10'd32;    
		mem[   412] = 10'd33;    
		mem[   413] = 10'd32;    
		mem[   414] = 10'd33;    
		mem[   415] = 10'd32;    
		mem[   416] = 10'd33;    
		mem[   417] = 10'd32;    
		mem[   418] = 10'd33;    
		mem[   419] = 10'd32;    
		mem[   420] = 10'd33;    
		mem[   421] = 10'd32;    
		mem[   422] = 10'd32;    
		mem[   423] = 10'd33;    
		mem[   424] = 10'd33;    
		mem[   425] = 10'd32;    
		mem[   426] = 10'd33;    
		mem[   427] = 10'd32;    
		mem[   428] = 10'd32;    
		mem[   429] = 10'd33;    
		mem[   430] = 10'd32;    
		mem[   431] = 10'd33;    
		mem[   432] = 10'd32;    
		mem[   433] = 10'd33;    
		mem[   434] = 10'd32;    
		mem[   435] = 10'd33;    
		mem[   436] = 10'd32;    
		mem[   437] = 10'd33;    
		mem[   438] = 10'd32;    
		mem[   439] = 10'd33;    
		mem[   440] = 10'd32;    
		mem[   441] = 10'd33;    
		mem[   442] = 10'd32;    
		mem[   443] = 10'd33;    
		mem[   444] = 10'd32;    
		mem[   445] = 10'd33;    
		mem[   446] = 10'd32;    
		mem[   447] = 10'd33;    
		mem[   448] = 10'd32;    
		mem[   449] = 10'd33;    
		mem[   450] = 10'd32;    
		mem[   451] = 10'd33;    
		mem[   452] = 10'd32;    
		mem[   453] = 10'd33;    
		mem[   454] = 10'd32;    
		mem[   455] = 10'd33;    
		mem[   456] = 10'd32;    
		mem[   457] = 10'd70;    
		mem[   458] = 10'd28;    
		mem[   459] = 10'd107;    
		mem[   460] = 10'd83;    
		mem[   461] = 10'd27;    
		mem[   462] = 10'd108;    
		mem[   463] = 10'd83;    
		mem[   464] = 10'd28;    
		mem[   465] = 10'd108;    
		mem[   466] = 10'd83;    
		mem[   467] = 10'd27;    
		mem[   468] = 10'd109;    
		mem[   469] = 10'd82;    
		mem[   470] = 10'd28;    
		mem[   471] = 10'd108;    
		mem[   472] = 10'd83;    
		mem[   473] = 10'd28;    
		mem[   474] = 10'd108;    
		mem[   475] = 10'd82;    
		mem[   476] = 10'd28;    
		mem[   477] = 10'd108;    
		mem[   478] = 10'd83;    
		mem[   479] = 10'd28;    
		mem[   480] = 10'd108;    
		mem[   481] = 10'd82;    
		mem[   482] = 10'd27;    
		mem[   483] = 10'd109;    
		mem[   484] = 10'd83;    
		mem[   485] = 10'd27;    
		mem[   486] = 10'd109;    
		mem[   487] = 10'd82;    
		mem[   488] = 10'd28;    
		mem[   489] = 10'd108;    
		mem[   490] = 10'd83;    
		mem[   491] = 10'd27;    
		mem[   492] = 10'd108;    
		mem[   493] = 10'd83;    
		mem[   494] = 10'd28;    
		mem[   495] = 10'd108;    
		mem[   496] = 10'd83;    
		mem[   497] = 10'd41;    
		mem[   498] = 10'd36;    
		mem[   499] = 10'd47;    
		mem[   500] = 10'd38;    
		mem[   501] = 10'd32;    
		mem[   502] = 10'd36;    
		mem[   503] = 10'd49;    
		mem[   504] = 10'd31;    
		mem[   505] = 10'd39;    
		mem[   506] = 10'd82;    
		mem[   507] = 10'd40;    
		mem[   508] = 10'd33;    
		mem[   509] = 10'd36;    
		mem[   510] = 10'd49;    
		mem[   511] = 10'd31;    
		mem[   512] = 10'd40;    
		mem[   513] = 10'd35;    
		mem[   514] = 10'd48;    
		mem[   515] = 10'd39;    
		mem[   516] = 10'd33;    
		mem[   517] = 10'd37;    
		mem[   518] = 10'd48;    
		mem[   519] = 10'd31;    
		mem[   520] = 10'd40;    
		mem[   521] = 10'd35;    
		mem[   522] = 10'd48;    
		mem[   523] = 10'd39;    
		mem[   524] = 10'd33;    
		mem[   525] = 10'd37;    
		mem[   526] = 10'd47;    
		mem[   527] = 10'd32;    
		mem[   528] = 10'd40;    
		mem[   529] = 10'd36;    
		mem[   530] = 10'd46;    
		mem[   531] = 10'd40;    
		mem[   532] = 10'd33;    
		mem[   533] = 10'd37;    
		mem[   534] = 10'd74;    
		mem[   535] = 10'd40;    
		mem[   536] = 10'd150;    
		mem[   537] = 10'd117;    
		mem[   538] = 10'd39;    
		mem[   539] = 10'd154;    
		mem[   540] = 10'd118;    
		mem[   541] = 10'd39;    
		mem[   542] = 10'd155;    
		mem[   543] = 10'd117;    
		mem[   544] = 10'd39;    
		mem[   545] = 10'd154;    
		mem[   546] = 10'd118;    
		mem[   547] = 10'd39;    
		mem[   548] = 10'd107;    
		mem[   549] = 10'd19;    
		mem[   550] = 10'd19;    
		mem[   551] = 10'd19;    
		mem[   552] = 10'd18;    
		mem[   553] = 10'd20;    
		mem[   554] = 10'd21;    
		mem[   555] = 10'd20;    
		mem[   556] = 10'd19;    
		mem[   557] = 10'd18;    
		mem[   558] = 10'd21;    
		mem[   559] = 10'd18;    
		mem[   560] = 10'd19;    
		mem[   561] = 10'd19;    
		mem[   562] = 10'd20;    
		mem[   563] = 10'd21;    
		mem[   564] = 10'd20;    
		mem[   565] = 10'd19;    
		mem[   566] = 10'd18;    
		mem[   567] = 10'd19;    
		mem[   568] = 10'd19;    
		mem[   569] = 10'd19;    
		mem[   570] = 10'd21;    
		mem[   571] = 10'd19;    
		mem[   572] = 10'd19;    
		mem[   573] = 10'd19;    
		mem[   574] = 10'd20;    
		mem[   575] = 10'd19;    
		mem[   576] = 10'd18;    
		mem[   577] = 10'd20;    
		mem[   578] = 10'd19;    
		mem[   579] = 10'd20;    
		mem[   580] = 10'd20;    
		mem[   581] = 10'd20;    
		mem[   582] = 10'd19;    
		mem[   583] = 10'd18;    
		mem[   584] = 10'd19;    
		mem[   585] = 10'd19;    
		mem[   586] = 10'd20;    
		mem[   587] = 10'd20;    
		mem[   588] = 10'd20;    
		mem[   589] = 10'd18;    
		mem[   590] = 10'd20;    
		mem[   591] = 10'd19;    
		mem[   592] = 10'd19;    
		mem[   593] = 10'd19;    
		mem[   594] = 10'd20;    
		mem[   595] = 10'd20;    
		mem[   596] = 10'd19;    
		mem[   597] = 10'd20;    
		mem[   598] = 10'd19;    
		mem[   599] = 10'd18;    
		mem[   600] = 10'd19;    
		mem[   601] = 10'd20;    
		mem[   602] = 10'd20;    
		mem[   603] = 10'd20;    
		mem[   604] = 10'd19;    
		mem[   605] = 10'd18;    
		mem[   606] = 10'd20;    
		mem[   607] = 10'd19;    
		mem[   608] = 10'd19;    
		mem[   609] = 10'd19;    
		mem[   610] = 10'd20;    
		mem[   611] = 10'd20;    
		mem[   612] = 10'd19;    
		mem[   613] = 10'd20;    
		mem[   614] = 10'd19;    
		mem[   615] = 10'd19;    
		mem[   616] = 10'd18;    
		mem[   617] = 10'd20;    
		mem[   618] = 10'd20;    
		mem[   619] = 10'd20;    
		mem[   620] = 10'd19;    
		mem[   621] = 10'd19;    
		mem[   622] = 10'd19;    
		mem[   623] = 10'd19;    
		mem[   624] = 10'd279;    
		mem[   625] = 10'd878;    
		mem[   626] = 10'd354;    
		mem[   627] = 10'd24;    
		mem[   628] = 10'd25;    
		mem[   629] = 10'd25;    
		mem[   630] = 10'd25;    
		mem[   631] = 10'd26;    
		mem[   632] = 10'd25;    
		mem[   633] = 10'd26;    
		mem[   634] = 10'd25;    
		mem[   635] = 10'd26;    
		mem[   636] = 10'd26;    
		mem[   637] = 10'd26;    
		mem[   638] = 10'd25;    
		mem[   639] = 10'd26;    
		mem[   640] = 10'd26;    
		mem[   641] = 10'd26;    
		mem[   642] = 10'd26;    
		mem[   643] = 10'd25;    
		mem[   644] = 10'd26;    
		mem[   645] = 10'd26;    
		mem[   646] = 10'd26;    
		mem[   647] = 10'd26;    
		mem[   648] = 10'd26;    
		mem[   649] = 10'd26;    
		mem[   650] = 10'd25;    
		mem[   651] = 10'd26;    
		mem[   652] = 10'd26;    
		mem[   653] = 10'd26;    
		mem[   654] = 10'd26;    
		mem[   655] = 10'd25;    
		mem[   656] = 10'd26;    
		mem[   657] = 10'd26;    
		mem[   658] = 10'd26;    
		mem[   659] = 10'd26;    
		mem[   660] = 10'd26;    
		mem[   661] = 10'd26;    
		mem[   662] = 10'd25;    
		mem[   663] = 10'd26;    
		mem[   664] = 10'd26;    
		mem[   665] = 10'd26;    
		mem[   666] = 10'd26;    
		mem[   667] = 10'd26;    
		mem[   668] = 10'd25;    
		mem[   669] = 10'd26;    
		mem[   670] = 10'd26;    
		mem[   671] = 10'd26;    
		mem[   672] = 10'd26;    
		mem[   673] = 10'd25;    
		mem[   674] = 10'd26;    
		mem[   675] = 10'd26;    
		mem[   676] = 10'd26;    
		mem[   677] = 10'd26;    
		mem[   678] = 10'd26;    
		mem[   679] = 10'd25;    
		mem[   680] = 10'd26;    
		mem[   681] = 10'd211;    
		mem[   682] = 10'd1023;//10'd1272;    
		mem[   683] = 10'd28;    
		mem[   684] = 10'd30;    
		mem[   685] = 10'd69;    
		mem[   686] = 10'd27;    
		mem[   687] = 10'd66;    
		mem[   688] = 10'd21;    
		mem[   689] = 10'd32;    
		mem[   690] = 10'd34;    
		mem[   691] = 10'd36;    
		mem[   692] = 10'd25;    
		mem[   693] = 10'd30;    
		mem[   694] = 10'd35;    
		mem[   695] = 10'd31;    
		mem[   696] = 10'd23;    
		mem[   697] = 10'd37;    
		mem[   698] = 10'd32;    
		mem[   699] = 10'd24;    
		mem[   700] = 10'd37;    
		mem[   701] = 10'd29;    
		mem[   702] = 10'd29;    
		mem[   703] = 10'd26;    
		mem[   704] = 10'd39;    
		mem[   705] = 10'd29;    
		mem[   706] = 10'd24;    
		mem[   707] = 10'd39;    
		mem[   708] = 10'd26;    
		mem[   709] = 10'd30;    
		mem[   710] = 10'd30;    
		mem[   711] = 10'd37;    
		mem[   712] = 10'd27;    
		mem[   713] = 10'd26;    
		mem[   714] = 10'd38;    
		mem[   715] = 10'd22;    
		mem[   716] = 10'd33;    
		mem[   717] = 10'd33;    
		mem[   718] = 10'd35;    
		mem[   719] = 10'd25;    
		mem[   720] = 10'd31;    
		mem[   721] = 10'd34;    
		mem[   722] = 10'd31;    
		mem[   723] = 10'd25;    
		mem[   724] = 10'd36;    
		mem[   725] = 10'd31;    
		mem[   726] = 10'd25;    
		mem[   727] = 10'd36;    
		mem[   728] = 10'd54;    
		mem[   729] = 10'd104;    
		mem[   730] = 10'd79;    
		mem[   731] = 10'd29;    
		mem[   732] = 10'd103;    
		mem[   733] = 10'd78;    
		mem[   734] = 10'd26;    
		mem[   735] = 10'd103;    
		mem[   736] = 10'd77;    
		mem[   737] = 10'd26;    
		mem[   738] = 10'd100;    
		mem[   739] = 10'd77;    
		mem[   740] = 10'd27;    
		mem[   741] = 10'd102;    
		mem[   742] = 10'd77;    
		mem[   743] = 10'd27;    
		mem[   744] = 10'd102;    
		mem[   745] = 10'd78;    
		mem[   746] = 10'd29;    
		mem[   747] = 10'd100;    
		mem[   748] = 10'd84;    
		mem[   749] = 10'd18;    
		mem[   750] = 10'd19;    
		mem[   751] = 10'd17;    
		mem[   752] = 10'd19;    
		mem[   753] = 10'd19;    
		mem[   754] = 10'd22;    
		mem[   755] = 10'd22;    
		mem[   756] = 10'd36;    
		mem[   757] = 10'd18;    
		mem[   758] = 10'd17;    
		mem[   759] = 10'd39;    
		mem[   760] = 10'd24;    
		mem[   761] = 10'd19;    
		mem[   762] = 10'd17;    
		mem[   763] = 10'd40;    
		mem[   764] = 10'd15;    
		mem[   765] = 10'd39;    
		mem[   766] = 10'd21;    
		mem[   767] = 10'd22;    
		mem[   768] = 10'd20;    
		mem[   769] = 10'd18;    
		mem[   770] = 10'd18;    
		mem[   771] = 10'd16;    
		mem[   772] = 10'd41;    
		mem[   773] = 10'd22;    
		mem[   774] = 10'd20;    
		mem[   775] = 10'd18;    
		mem[   776] = 10'd12;    
		mem[   777] = 10'd27;    
		mem[   778] = 10'd16;    
		mem[   779] = 10'd38;    
		mem[   780] = 10'd21;    
		mem[   781] = 10'd22;    
		mem[   782] = 10'd20;    
		mem[   783] = 10'd19;    
		mem[   784] = 10'd18;    
		mem[   785] = 10'd16;    
		mem[   786] = 10'd40;    
		mem[   787] = 10'd22;    
		mem[   788] = 10'd20;    
		mem[   789] = 10'd18;    
		mem[   790] = 10'd15;    
		mem[   791] = 10'd25;    
		mem[   792] = 10'd16;    
		mem[   793] = 10'd18;    
		mem[   794] = 10'd20;    
		mem[   795] = 10'd21;    
		mem[   796] = 10'd21;    
		mem[   797] = 10'd20;    
		mem[   798] = 10'd19;    
		mem[   799] = 10'd18;    
		mem[   800] = 10'd17;    
		mem[   801] = 10'd18;    
		mem[   802] = 10'd21;    
		mem[   803] = 10'd22;    
		mem[   804] = 10'd20;    
		mem[   805] = 10'd18;    
		mem[   806] = 10'd16;    
		mem[   807] = 10'd24;    
		mem[   808] = 10'd16;    
		mem[   809] = 10'd18;    
		mem[   810] = 10'd20;    
		mem[   811] = 10'd21;    
		mem[   812] = 10'd21;    
		mem[   813] = 10'd20;    
		mem[   814] = 10'd19;    
		mem[   815] = 10'd18;    
		mem[   816] = 10'd18;    
		mem[   817] = 10'd25;    
		mem[   818] = 10'd29;    
		mem[   819] = 10'd29;    
		mem[   820] = 10'd23;    
		mem[   821] = 10'd25;    
		mem[   822] = 10'd25;    
		mem[   823] = 10'd24;    
		mem[   824] = 10'd28;    
		mem[   825] = 10'd28;    
		mem[   826] = 10'd28;    
		mem[   827] = 10'd24;    
		mem[   828] = 10'd22;    
		mem[   829] = 10'd24;    
		mem[   830] = 10'd30;    
		mem[   831] = 10'd28;    
		mem[   832] = 10'd24;    
		mem[   833] = 10'd25;    
		mem[   834] = 10'd25;    
		mem[   835] = 10'd24;    
		mem[   836] = 10'd27;    
		mem[   837] = 10'd29;    
		mem[   838] = 10'd27;    
		mem[   839] = 10'd24;    
		mem[   840] = 10'd23;    
		mem[   841] = 10'd25;    
		mem[   842] = 10'd29;    
		mem[   843] = 10'd28;    
		mem[   844] = 10'd24;    
		mem[   845] = 10'd24;    
		mem[   846] = 10'd26;    
		mem[   847] = 10'd24;    
		mem[   848] = 10'd27;    
		mem[   849] = 10'd28;    
		mem[   850] = 10'd27;    
		mem[   851] = 10'd25;    
		mem[   852] = 10'd23;    
		mem[   853] = 10'd25;    
		mem[   854] = 10'd29;    
		mem[   855] = 10'd27;    
		mem[   856] = 10'd25;    
		mem[   857] = 10'd24;    
		mem[   858] = 10'd26;    
		mem[   859] = 10'd24;    
		mem[   860] = 10'd27;    
		mem[   861] = 10'd28;    
		mem[   862] = 10'd26;    
		mem[   863] = 10'd25;    
		mem[   864] = 10'd25;    
		mem[   865] = 10'd24;    
		mem[   866] = 10'd28;    
		mem[   867] = 10'd27;    
		mem[   868] = 10'd25;    
		mem[   869] = 10'd25;    
		mem[   870] = 10'd26;    
		mem[   871] = 10'd24;    
		mem[   872] = 10'd27;    
		mem[   873] = 10'd213;    
		mem[   874] = 10'd47;    
		mem[   875] = 10'd156;    
		mem[   876] = 10'd116;    
		mem[   877] = 10'd39;    
		mem[   878] = 10'd154;    
		mem[   879] = 10'd112;    
		mem[   880] = 10'd40;    
		mem[   881] = 10'd152;    
		mem[   882] = 10'd116;    
		mem[   883] = 10'd42;    
		mem[   884] = 10'd154;    
		mem[   885] = 10'd115;    
		mem[   886] = 10'd39;    
		mem[   887] = 10'd154;    
		mem[   888] = 10'd120;    
		mem[   889] = 10'd38;    
		mem[   890] = 10'd1023;//10'd1141;    
		mem[   891] = 10'd29;    
		mem[   892] = 10'd30;    
		mem[   893] = 10'd30;    
		mem[   894] = 10'd30;    
		mem[   895] = 10'd30;    
		mem[   896] = 10'd31;    
		mem[   897] = 10'd30;    
		mem[   898] = 10'd31;    
		mem[   899] = 10'd30;    
		mem[   900] = 10'd31;    
		mem[   901] = 10'd30;    
		mem[   902] = 10'd31;    
		mem[   903] = 10'd31;    
		mem[   904] = 10'd31;    
		mem[   905] = 10'd30;    
		mem[   906] = 10'd31;    
		mem[   907] = 10'd30;    
		mem[   908] = 10'd31;    
		mem[   909] = 10'd31;    
		mem[   910] = 10'd30;    
		mem[   911] = 10'd31;    
		mem[   912] = 10'd31;    
		mem[   913] = 10'd30;    
		mem[   914] = 10'd31;    
		mem[   915] = 10'd31;    
		mem[   916] = 10'd30;    
		mem[   917] = 10'd31;    
		mem[   918] = 10'd31;    
		mem[   919] = 10'd30;    
		mem[   920] = 10'd31;    
		mem[   921] = 10'd31;    
		mem[   922] = 10'd30;    
		mem[   923] = 10'd31;    
		mem[   924] = 10'd31;    
		mem[   925] = 10'd30;    
		mem[   926] = 10'd31;    
		mem[   927] = 10'd31;    
		mem[   928] = 10'd30;    
		mem[   929] = 10'd31;    
		mem[   930] = 10'd30;    
		mem[   931] = 10'd31;    
		mem[   932] = 10'd31;    
		mem[   933] = 10'd30;    
		mem[   934] = 10'd31;    
		mem[   935] = 10'd31;    
		mem[   936] = 10'd30;    
		mem[   937] = 10'd31;    
		mem[   938] = 10'd31;    
		mem[   939] = 10'd30;    
		mem[   940] = 10'd31;    
		mem[   941] = 10'd31;    
		mem[   942] = 10'd30;    
		mem[   943] = 10'd31;    
		mem[   944] = 10'd30;    
		mem[   945] = 10'd31;    
		mem[   946] = 10'd31;    
		mem[   947] = 10'd30;    
		mem[   948] = 10'd31;    
		mem[   949] = 10'd31;    
		mem[   950] = 10'd30;    
		mem[   951] = 10'd31;    
		mem[   952] = 10'd31;    
		mem[   953] = 10'd30;    
		mem[   954] = 10'd31;    
		mem[   955] = 10'd30;    
		mem[   956] = 10'd31;    
		mem[   957] = 10'd31;    
		mem[   958] = 10'd30;    
		mem[   959] = 10'd31;    
		mem[   960] = 10'd31;    
		mem[   961] = 10'd30;    
		mem[   962] = 10'd31;    
		mem[   963] = 10'd31;    
		mem[   964] = 10'd30;    
		mem[   965] = 10'd31;    
		mem[   966] = 10'd30;    
		mem[   967] = 10'd31;    
		mem[   968] = 10'd31;    
		mem[   969] = 10'd30;    
		mem[   970] = 10'd31;    
		mem[   971] = 10'd31;    
		mem[   972] = 10'd30;    
		mem[   973] = 10'd31;    
		mem[   974] = 10'd31;    
		mem[   975] = 10'd30;    
		mem[   976] = 10'd31;    
		mem[   977] = 10'd31;    
		mem[   978] = 10'd30;    
		mem[   979] = 10'd31;    
		mem[   980] = 10'd30;    
		mem[   981] = 10'd31;    
		mem[   982] = 10'd31;    
		mem[   983] = 10'd30;    
		mem[   984] = 10'd31;    
		mem[   985] = 10'd70;    
		mem[   986] = 10'd27;    
		mem[   987] = 10'd102;    
		mem[   988] = 10'd78;    
		mem[   989] = 10'd27;    
		mem[   990] = 10'd101;    
		mem[   991] = 10'd78;    
		mem[   992] = 10'd27;    
		mem[   993] = 10'd102;    
		mem[   994] = 10'd78;    
		mem[   995] = 10'd26;    
		mem[   996] = 10'd102;    
		mem[   997] = 10'd79;    
		mem[   998] = 10'd26;    
		mem[   999] = 10'd102;    
		mem[  1000] = 10'd78;    
		mem[  1001] = 10'd26;    
		mem[  1002] = 10'd102;    
		mem[  1003] = 10'd78;    
		mem[  1004] = 10'd26;    
		mem[  1005] = 10'd103;    
		mem[  1006] = 10'd78;    
		mem[  1007] = 10'd26;    
		mem[  1008] = 10'd103;    
		mem[  1009] = 10'd77;    
		mem[  1010] = 10'd27;    
		mem[  1011] = 10'd102;    
		mem[  1012] = 10'd78;    
		mem[  1013] = 10'd26;    
		mem[  1014] = 10'd102;    
		mem[  1015] = 10'd78;    
		mem[  1016] = 10'd27;    
		mem[  1017] = 10'd102;    
		mem[  1018] = 10'd78;    
		mem[  1019] = 10'd26;    
		mem[  1020] = 10'd102;    
		mem[  1021] = 10'd78;    
		mem[  1022] = 10'd26;    
		mem[  1023] = 10'd103;    
		mem[  1024] = 10'd78;    
		mem[  1025] = 10'd26;    
		mem[  1026] = 10'd103;    
		mem[  1027] = 10'd107;    
		mem[  1028] = 10'd41;    
		mem[  1029] = 10'd37;    
		mem[  1030] = 10'd50;    
		mem[  1031] = 10'd41;    
		mem[  1032] = 10'd35;    
		mem[  1033] = 10'd89;    
		mem[  1034] = 10'd33;    
		mem[  1035] = 10'd42;    
		mem[  1036] = 10'd87;    
		mem[  1037] = 10'd41;    
		mem[  1038] = 10'd35;    
		mem[  1039] = 10'd38;    
		mem[  1040] = 10'd52;    
		mem[  1041] = 10'd33;    
		mem[  1042] = 10'd42;    
		mem[  1043] = 10'd36;    
		mem[  1044] = 10'd50;    
		mem[  1045] = 10'd42;    
		mem[  1046] = 10'd35;    
		mem[  1047] = 10'd39;    
		mem[  1048] = 10'd50;    
		mem[  1049] = 10'd34;    
		mem[  1050] = 10'd42;    
		mem[  1051] = 10'd37;    
		mem[  1052] = 10'd49;    
		mem[  1053] = 10'd41;    
		mem[  1054] = 10'd36;    
		mem[  1055] = 10'd39;    
		mem[  1056] = 10'd49;    
		mem[  1057] = 10'd35;    
		mem[  1058] = 10'd41;    
		mem[  1059] = 10'd38;    
		mem[  1060] = 10'd117;    
		mem[  1061] = 10'd122;    
		mem[  1062] = 10'd42;    
		mem[  1063] = 10'd162;    
		mem[  1064] = 10'd124;    
		mem[  1065] = 10'd41;    
		mem[  1066] = 10'd163;    
		mem[  1067] = 10'd124;    
		mem[  1068] = 10'd42;    
		mem[  1069] = 10'd161;    
		mem[  1070] = 10'd124;    
		mem[  1071] = 10'd42;    
		mem[  1072] = 10'd163;    
		mem[  1073] = 10'd53;    
		mem[  1074] = 10'd22;    
		mem[  1075] = 10'd21;    
		mem[  1076] = 10'd20;    
		mem[  1077] = 10'd19;    
		mem[  1078] = 10'd23;    
		mem[  1079] = 10'd19;    
		mem[  1080] = 10'd20;    
		mem[  1081] = 10'd21;    
		mem[  1082] = 10'd21;    
		mem[  1083] = 10'd21;    
		mem[  1084] = 10'd21;    
		mem[  1085] = 10'd20;    
		mem[  1086] = 10'd20;    
		mem[  1087] = 10'd20;    
		mem[  1088] = 10'd20;    
		mem[  1089] = 10'd21;    
		mem[  1090] = 10'd22;    
		mem[  1091] = 10'd20;    
		mem[  1092] = 10'd20;    
		mem[  1093] = 10'd19;    
		mem[  1094] = 10'd23;    
		mem[  1095] = 10'd19;    
		mem[  1096] = 10'd20;    
		mem[  1097] = 10'd21;    
		mem[  1098] = 10'd21;    
		mem[  1099] = 10'd21;    
		mem[  1100] = 10'd21;    
		mem[  1101] = 10'd20;    
		mem[  1102] = 10'd20;    
		mem[  1103] = 10'd19;    
		mem[  1104] = 10'd20;    
		mem[  1105] = 10'd22;    
		mem[  1106] = 10'd21;    
		mem[  1107] = 10'd21;    
		mem[  1108] = 10'd20;    
		mem[  1109] = 10'd19;    
		mem[  1110] = 10'd22;    
		mem[  1111] = 10'd19;    
		mem[  1112] = 10'd21;    
		mem[  1113] = 10'd20;    
		mem[  1114] = 10'd21;    
		mem[  1115] = 10'd21;    
		mem[  1116] = 10'd21;    
		mem[  1117] = 10'd20;    
		mem[  1118] = 10'd20;    
		mem[  1119] = 10'd20;    
		mem[  1120] = 10'd20;    
		mem[  1121] = 10'd21;    
		mem[  1122] = 10'd22;    
		mem[  1123] = 10'd20;    
		mem[  1124] = 10'd20;    
		mem[  1125] = 10'd20;    
		mem[  1126] = 10'd22;    
		mem[  1127] = 10'd19;    
		mem[  1128] = 10'd20;    
		mem[  1129] = 10'd21;    
		mem[  1130] = 10'd21;    
		mem[  1131] = 10'd21;    
		mem[  1132] = 10'd20;    
		mem[  1133] = 10'd21;    
		mem[  1134] = 10'd20;    
		mem[  1135] = 10'd20;    
		mem[  1136] = 10'd20;    
		mem[  1137] = 10'd21;    
		mem[  1138] = 10'd21;    
		mem[  1139] = 10'd21;    
		mem[  1140] = 10'd20;    
		mem[  1141] = 10'd20;    
		mem[  1142] = 10'd21;    
		mem[  1143] = 10'd20;    
		mem[  1144] = 10'd282;    
		mem[  1145] = 10'd44;    
		mem[  1146] = 10'd174;    
		mem[  1147] = 10'd112;    
		mem[  1148] = 10'd42;    
		mem[  1149] = 10'd861;    
		mem[  1150] = 10'd26;    
		mem[  1151] = 10'd26;    
		mem[  1152] = 10'd27;    
		mem[  1153] = 10'd27;    
		mem[  1154] = 10'd27;    
		mem[  1155] = 10'd27;    
		mem[  1156] = 10'd27;    
		mem[  1157] = 10'd27;    
		mem[  1158] = 10'd27;    
		mem[  1159] = 10'd27;    
		mem[  1160] = 10'd27;    
		mem[  1161] = 10'd28;    
		mem[  1162] = 10'd27;    
		mem[  1163] = 10'd27;    
		mem[  1164] = 10'd28;    
		mem[  1165] = 10'd27;    
		mem[  1166] = 10'd27;    
		mem[  1167] = 10'd28;    
		mem[  1168] = 10'd27;    
		mem[  1169] = 10'd27;    
		mem[  1170] = 10'd28;    
		mem[  1171] = 10'd27;    
		mem[  1172] = 10'd27;    
		mem[  1173] = 10'd28;    
		mem[  1174] = 10'd27;    
		mem[  1175] = 10'd28;    
		mem[  1176] = 10'd27;    
		mem[  1177] = 10'd27;    
		mem[  1178] = 10'd27;    
		mem[  1179] = 10'd28;    
		mem[  1180] = 10'd27;    
		mem[  1181] = 10'd27;    
		mem[  1182] = 10'd28;    
		mem[  1183] = 10'd27;    
		mem[  1184] = 10'd27;    
		mem[  1185] = 10'd28;    
		mem[  1186] = 10'd27;    
		mem[  1187] = 10'd28;    
		mem[  1188] = 10'd27;    
		mem[  1189] = 10'd27;    
		mem[  1190] = 10'd27;    
		mem[  1191] = 10'd28;    
		mem[  1192] = 10'd27;    
		mem[  1193] = 10'd27;    
		mem[  1194] = 10'd28;    
		mem[  1195] = 10'd27;    
		mem[  1196] = 10'd27;    
		mem[  1197] = 10'd28;    
		mem[  1198] = 10'd27;    
		mem[  1199] = 10'd27;    
		mem[  1200] = 10'd28;    
		mem[  1201] = 10'd1023;// 10'd1484;    
		mem[  1202] = 10'd69;    
		mem[  1203] = 10'd31;    
		mem[  1204] = 10'd27;    
		mem[  1205] = 10'd43;    
		mem[  1206] = 10'd29;    
		mem[  1207] = 10'd69;    
		mem[  1208] = 10'd25;    
		mem[  1209] = 10'd32;    
		mem[  1210] = 10'd32;    
		mem[  1211] = 10'd41;    
		mem[  1212] = 10'd26;    
		mem[  1213] = 10'd69;    
		mem[  1214] = 10'd21;    
		mem[  1215] = 10'd8;    
		mem[  1216] = 10'd29;    
		mem[  1217] = 10'd37;    
		mem[  1218] = 10'd36;    
		mem[  1219] = 10'd25;    
		mem[  1220] = 10'd36;    
		mem[  1221] = 10'd34;    
		mem[  1222] = 10'd32;    
		mem[  1223] = 10'd27;    
		mem[  1224] = 10'd39;    
		mem[  1225] = 10'd33;    
		mem[  1226] = 10'd25;    
		mem[  1227] = 10'd41;    
		mem[  1228] = 10'd28;    
		mem[  1229] = 10'd32;    
		mem[  1230] = 10'd30;    
		mem[  1231] = 10'd40;    
		mem[  1232] = 10'd29;    
		mem[  1233] = 10'd27;    
		mem[  1234] = 10'd42;    
		mem[  1235] = 10'd24;    
		mem[  1236] = 10'd34;    
		mem[  1237] = 10'd34;    
		mem[  1238] = 10'd38;    
		mem[  1239] = 10'd28;    
		mem[  1240] = 10'd31;    
		mem[  1241] = 10'd37;    
		mem[  1242] = 10'd33;    
		mem[  1243] = 10'd25;    
		mem[  1244] = 10'd79;    
		mem[  1245] = 10'd91;    
		mem[  1246] = 10'd28;    
		mem[  1247] = 10'd112;    
		mem[  1248] = 10'd80;    
		mem[  1249] = 10'd31;    
		mem[  1250] = 10'd108;    
		mem[  1251] = 10'd82;    
		mem[  1252] = 10'd28;    
		mem[  1253] = 10'd105;    
		mem[  1254] = 10'd82;    
		mem[  1255] = 10'd30;    
		mem[  1256] = 10'd106;    
		mem[  1257] = 10'd82;    
		mem[  1258] = 10'd28;    
		mem[  1259] = 10'd108;    
		mem[  1260] = 10'd82;    
		mem[  1261] = 10'd29;    
		mem[  1262] = 10'd108;    
		mem[  1263] = 10'd90;    
		mem[  1264] = 10'd20;    
		mem[  1265] = 10'd20;    
		mem[  1266] = 10'd17;    
		mem[  1267] = 10'd20;    
		mem[  1268] = 10'd21;    
		mem[  1269] = 10'd23;    
		mem[  1270] = 10'd23;    
		mem[  1271] = 10'd21;    
		mem[  1272] = 10'd18;    
		mem[  1273] = 10'd18;    
		mem[  1274] = 10'd18;    
		mem[  1275] = 10'd44;    
		mem[  1276] = 10'd23;    
		mem[  1277] = 10'd20;    
		mem[  1278] = 10'd18;    
		mem[  1279] = 10'd41;    
		mem[  1280] = 10'd18;    
		mem[  1281] = 10'd41;    
		mem[  1282] = 10'd24;    
		mem[  1283] = 10'd22;    
		mem[  1284] = 10'd21;    
		mem[  1285] = 10'd19;    
		mem[  1286] = 10'd18;    
		mem[  1287] = 10'd18;    
		mem[  1288] = 10'd45;    
		mem[  1289] = 10'd23;    
		mem[  1290] = 10'd19;    
		mem[  1291] = 10'd18;    
		mem[  1292] = 10'd42;    
		mem[  1293] = 10'd18;    
		mem[  1294] = 10'd20;    
		mem[  1295] = 10'd21;    
		mem[  1296] = 10'd23;    
		mem[  1297] = 10'd23;    
		mem[  1298] = 10'd21;    
		mem[  1299] = 10'd19;    
		mem[  1300] = 10'd18;    
		mem[  1301] = 10'd19;    
		mem[  1302] = 10'd43;    
		mem[  1303] = 10'd23;    
		mem[  1304] = 10'd20;    
		mem[  1305] = 10'd18;    
		mem[  1306] = 10'd41;    
		mem[  1307] = 10'd19;    
		mem[  1308] = 10'd20;    
		mem[  1309] = 10'd21;    
		mem[  1310] = 10'd23;    
		mem[  1311] = 10'd22;    
		mem[  1312] = 10'd21;    
		mem[  1313] = 10'd19;    
		mem[  1314] = 10'd19;    
		mem[  1315] = 10'd19;    
		mem[  1316] = 10'd19;    
		mem[  1317] = 10'd24;    
		mem[  1318] = 10'd23;    
		mem[  1319] = 10'd20;    
		mem[  1320] = 10'd18;    
		mem[  1321] = 10'd41;    
		mem[  1322] = 10'd19;    
		mem[  1323] = 10'd20;    
		mem[  1324] = 10'd21;    
		mem[  1325] = 10'd23;    
		mem[  1326] = 10'd26;    
		mem[  1327] = 10'd27;    
		mem[  1328] = 10'd25;    
		mem[  1329] = 10'd24;    
		mem[  1330] = 10'd29;    
		mem[  1331] = 10'd32;    
		mem[  1332] = 10'd26;    
		mem[  1333] = 10'd23;    
		mem[  1334] = 10'd31;    
		mem[  1335] = 10'd23;    
		mem[  1336] = 10'd28;    
		mem[  1337] = 10'd29;    
		mem[  1338] = 10'd30;    
		mem[  1339] = 10'd27;    
		mem[  1340] = 10'd26;    
		mem[  1341] = 10'd24;    
		mem[  1342] = 10'd29;    
		mem[  1343] = 10'd31;    
		mem[  1344] = 10'd26;    
		mem[  1345] = 10'd24;    
		mem[  1346] = 10'd30;    
		mem[  1347] = 10'd24;    
		mem[  1348] = 10'd28;    
		mem[  1349] = 10'd29;    
		mem[  1350] = 10'd30;    
		mem[  1351] = 10'd27;    
		mem[  1352] = 10'd25;    
		mem[  1353] = 10'd25;    
		mem[  1354] = 10'd28;    
		mem[  1355] = 10'd31;    
		mem[  1356] = 10'd27;    
		mem[  1357] = 10'd24;    
		mem[  1358] = 10'd30;    
		mem[  1359] = 10'd24;    
		mem[  1360] = 10'd27;    
		mem[  1361] = 10'd30;    
		mem[  1362] = 10'd29;    
		mem[  1363] = 10'd27;    
		mem[  1364] = 10'd26;    
		mem[  1365] = 10'd24;    
		mem[  1366] = 10'd29;    
		mem[  1367] = 10'd30;    
		mem[  1368] = 10'd27;    
		mem[  1369] = 10'd25;    
		mem[  1370] = 10'd30;    
		mem[  1371] = 10'd24;    
		mem[  1372] = 10'd28;    
		mem[  1373] = 10'd28;    
		mem[  1374] = 10'd30;    
		mem[  1375] = 10'd27;    
		mem[  1376] = 10'd26;    
		mem[  1377] = 10'd25;    
		mem[  1378] = 10'd28;    
		mem[  1379] = 10'd83;    
		mem[  1380] = 10'd48;    
		mem[  1381] = 10'd141;    
		mem[  1382] = 10'd118;    
		mem[  1383] = 10'd50;    
		mem[  1384] = 10'd154;    
		mem[  1385] = 10'd132;    
		mem[  1386] = 10'd42;    
		mem[  1387] = 10'd162;    
		mem[  1388] = 10'd124;    
		mem[  1389] = 10'd42;    
		mem[  1390] = 10'd162;    
		mem[  1391] = 10'd124;    
		mem[  1392] = 10'd42;    
		mem[  1393] = 10'd164;    
		mem[  1394] = 10'd122;    
		mem[  1395] = 10'd44;    
		mem[  1396] = 10'd1023;// 10'd1249;    
		mem[  1397] = 10'd35;    
		mem[  1398] = 10'd33;    
		mem[  1399] = 10'd34;    
		mem[  1400] = 10'd33;    
		mem[  1401] = 10'd32;    
		mem[  1402] = 10'd33;    
		mem[  1403] = 10'd33;    
		mem[  1404] = 10'd32;    
		mem[  1405] = 10'd33;    
		mem[  1406] = 10'd32;    
		mem[  1407] = 10'd33;    
		mem[  1408] = 10'd32;    
		mem[  1409] = 10'd33;    
		mem[  1410] = 10'd32;    
		mem[  1411] = 10'd33;    
		mem[  1412] = 10'd32;    
		mem[  1413] = 10'd32;    
		mem[  1414] = 10'd33;    
		mem[  1415] = 10'd32;    
		mem[  1416] = 10'd33;    
		mem[  1417] = 10'd32;    
		mem[  1418] = 10'd33;    
		mem[  1419] = 10'd32;    
		mem[  1420] = 10'd33;    
		mem[  1421] = 10'd32;    
		mem[  1422] = 10'd32;    
		mem[  1423] = 10'd33;    
		mem[  1424] = 10'd32;    
		mem[  1425] = 10'd33;    
		mem[  1426] = 10'd32;    
		mem[  1427] = 10'd33;    
		mem[  1428] = 10'd32;    
		mem[  1429] = 10'd33;    
		mem[  1430] = 10'd32;    
		mem[  1431] = 10'd33;    
		mem[  1432] = 10'd32;    
		mem[  1433] = 10'd33;    
		mem[  1434] = 10'd32;    
		mem[  1435] = 10'd32;    
		mem[  1436] = 10'd33;    
		mem[  1437] = 10'd32;    
		mem[  1438] = 10'd33;    
		mem[  1439] = 10'd32;    
		mem[  1440] = 10'd33;    
		mem[  1441] = 10'd32;    
		mem[  1442] = 10'd33;    
		mem[  1443] = 10'd32;    
		mem[  1444] = 10'd33;    
		mem[  1445] = 10'd32;    
		mem[  1446] = 10'd33;    
		mem[  1447] = 10'd32;    
		mem[  1448] = 10'd33;    
		mem[  1449] = 10'd32;    
		mem[  1450] = 10'd33;    
		mem[  1451] = 10'd32;    
		mem[  1452] = 10'd33;    
		mem[  1453] = 10'd32;    
		mem[  1454] = 10'd33;    
		mem[  1455] = 10'd32;    
		mem[  1456] = 10'd33;    
		mem[  1457] = 10'd32;    
		mem[  1458] = 10'd33;    
		mem[  1459] = 10'd32;    
		mem[  1460] = 10'd32;    
		mem[  1461] = 10'd33;    
		mem[  1462] = 10'd32;    
		mem[  1463] = 10'd33;    
		mem[  1464] = 10'd32;    
		mem[  1465] = 10'd33;    
		mem[  1466] = 10'd32;    
		mem[  1467] = 10'd33;    
		mem[  1468] = 10'd32;    
		mem[  1469] = 10'd33;    
		mem[  1470] = 10'd32;    
		mem[  1471] = 10'd33;    
		mem[  1472] = 10'd32;    
		mem[  1473] = 10'd33;    
		mem[  1474] = 10'd32;    
		mem[  1475] = 10'd33;    
		mem[  1476] = 10'd32;    
		mem[  1477] = 10'd33;    
		mem[  1478] = 10'd32;    
		mem[  1479] = 10'd33;    
		mem[  1480] = 10'd32;    
		mem[  1481] = 10'd33;    
		mem[  1482] = 10'd32;    
		mem[  1483] = 10'd33;    
		mem[  1484] = 10'd79;    
		mem[  1485] = 10'd28;    
		mem[  1486] = 10'd102;    
		mem[  1487] = 10'd82;    
		mem[  1488] = 10'd28;    
		mem[  1489] = 10'd107;    
		mem[  1490] = 10'd83;    
		mem[  1491] = 10'd28;    
		mem[  1492] = 10'd108;    
		mem[  1493] = 10'd83;    
		mem[  1494] = 10'd28;    
		mem[  1495] = 10'd108;    
		mem[  1496] = 10'd83;    
		mem[  1497] = 10'd28;    
		mem[  1498] = 10'd108;    
		mem[  1499] = 10'd82;    
		mem[  1500] = 10'd28;    
		mem[  1501] = 10'd109;    
		mem[  1502] = 10'd82;    
		mem[  1503] = 10'd28;    
		mem[  1504] = 10'd108;    
		mem[  1505] = 10'd83;    
		mem[  1506] = 10'd27;    
		mem[  1507] = 10'd109;    
		mem[  1508] = 10'd82;    
		mem[  1509] = 10'd28;    
		mem[  1510] = 10'd108;    
		mem[  1511] = 10'd83;    
		mem[  1512] = 10'd27;    
		mem[  1513] = 10'd109;    
		mem[  1514] = 10'd82;    
		mem[  1515] = 10'd27;    
		mem[  1516] = 10'd109;    
		mem[  1517] = 10'd82;    
		mem[  1518] = 10'd28;    
		mem[  1519] = 10'd108;    
		mem[  1520] = 10'd83;    
		mem[  1521] = 10'd30;    
		mem[  1522] = 10'd106;    
		mem[  1523] = 10'd83;    
		mem[  1524] = 10'd31;    
		mem[  1525] = 10'd76;    
		mem[  1526] = 10'd29;    
		mem[  1527] = 10'd31;    
		mem[  1528] = 10'd42;    
		mem[  1529] = 10'd34;    
		mem[  1530] = 10'd27;    
		mem[  1531] = 10'd45;    
		mem[  1532] = 10'd32;    
		mem[  1533] = 10'd26;    
		mem[  1534] = 10'd46;    
		mem[  1535] = 10'd24;    
		mem[  1536] = 10'd36;    
		mem[  1537] = 10'd39;    
		mem[  1538] = 10'd38;    
		mem[  1539] = 10'd27;    
		mem[  1540] = 10'd41;    
		mem[  1541] = 10'd31;    
		mem[  1542] = 10'd33;    
		mem[  1543] = 10'd34;    
		mem[  1544] = 10'd43;    
		mem[  1545] = 10'd28;    
		mem[  1546] = 10'd33;    
		mem[  1547] = 10'd39;    
		mem[  1548] = 10'd34;    
		mem[  1549] = 10'd28;    
		mem[  1550] = 10'd44;    
		mem[  1551] = 10'd32;    
		mem[  1552] = 10'd27;    
		mem[  1553] = 10'd45;    
		mem[  1554] = 10'd24;    
		mem[  1555] = 10'd37;    
		mem[  1556] = 10'd39;    
		mem[  1557] = 10'd37;    
		mem[  1558] = 10'd28;    
		mem[  1559] = 10'd41;    
		mem[  1560] = 10'd31;    
		mem[  1561] = 10'd33;    
		mem[  1562] = 10'd34;    
		mem[  1563] = 10'd42;    
		mem[  1564] = 10'd29;    
		mem[  1565] = 10'd33;    
		mem[  1566] = 10'd37;    
		mem[  1567] = 10'd32;    
		mem[  1568] = 10'd27;    
		mem[  1569] = 10'd37;    
		mem[  1570] = 10'd34;    
		mem[  1571] = 10'd27;    
		mem[  1572] = 10'd37;    
		mem[  1573] = 10'd31;    
		mem[  1574] = 10'd32;    
		mem[  1575] = 10'd29;    
		mem[  1576] = 10'd39;    
		mem[  1577] = 10'd31;    
		mem[  1578] = 10'd27;    
		mem[  1579] = 10'd39;    
		mem[  1580] = 10'd28;    
		mem[  1581] = 10'd33;    
		mem[  1582] = 10'd32;    
		mem[  1583] = 10'd38;    
		mem[  1584] = 10'd29;    
		mem[  1585] = 10'd30;    
		mem[  1586] = 10'd37;    
		mem[  1587] = 10'd30;    
		mem[  1588] = 10'd30;    
		mem[  1589] = 10'd35;    
		mem[  1590] = 10'd35;    
		mem[  1591] = 10'd28;    
		mem[  1592] = 10'd35;    
		mem[  1593] = 10'd34;    
		mem[  1594] = 10'd32;    
		mem[  1595] = 10'd28;    
		mem[  1596] = 10'd37;    
		mem[  1597] = 10'd33;    
		mem[  1598] = 10'd28;    
		mem[  1599] = 10'd36;    
		mem[  1600] = 10'd31;    
		mem[  1601] = 10'd32;    
		mem[  1602] = 10'd32;    
		mem[  1603] = 10'd36;    
		mem[  1604] = 10'd31;    
		mem[  1605] = 10'd30;    
		mem[  1606] = 10'd37;    
		mem[  1607] = 10'd28;    
		mem[  1608] = 10'd33;    
		mem[  1609] = 10'd33;    
		mem[  1610] = 10'd35;    
		mem[  1611] = 10'd28;    
		mem[  1612] = 10'd30;    
		mem[  1613] = 10'd33;    
		mem[  1614] = 10'd27;    
		mem[  1615] = 10'd32;    
		mem[  1616] = 10'd31;    
		mem[  1617] = 10'd33;    
		mem[  1618] = 10'd29;    
		mem[  1619] = 10'd29;    
		mem[  1620] = 10'd34;    
		mem[  1621] = 10'd28;    
		mem[  1622] = 10'd31;    
		mem[  1623] = 10'd30;    
		mem[  1624] = 10'd33;    
		mem[  1625] = 10'd30;    
		mem[  1626] = 10'd28;    
		mem[  1627] = 10'd34;    
		mem[  1628] = 10'd29;    
		mem[  1629] = 10'd30;    
		mem[  1630] = 10'd30;    
		mem[  1631] = 10'd33;    
		mem[  1632] = 10'd31;    
		mem[  1633] = 10'd28;    
		mem[  1634] = 10'd33;    
		mem[  1635] = 10'd30;    
		mem[  1636] = 10'd30;    
		mem[  1637] = 10'd30;    
		mem[  1638] = 10'd32;    
		mem[  1639] = 10'd31;    
		mem[  1640] = 10'd29;    
		mem[  1641] = 10'd32;    
		mem[  1642] = 10'd31;    
		mem[  1643] = 10'd30;    
		mem[  1644] = 10'd29;    
		mem[  1645] = 10'd32;    
		mem[  1646] = 10'd31;    
		mem[  1647] = 10'd30;    
		mem[  1648] = 10'd31;    
		mem[  1649] = 10'd31;    
		mem[  1650] = 10'd31;    
		mem[  1651] = 10'd29;    
		mem[  1652] = 10'd32;    
		mem[  1653] = 10'd31;    
		mem[  1654] = 10'd29;    
		mem[  1655] = 10'd31;    
		mem[  1656] = 10'd32;    
		mem[  1657] = 10'd30;    
		mem[  1658] = 10'd205;    
		mem[  1659] = 10'd31;    
		mem[  1660] = 10'd118;    
		mem[  1661] = 10'd838;    
		mem[  1662] = 10'd355;    
		mem[  1663] = 10'd34;    
		mem[  1664] = 10'd33;    
		mem[  1665] = 10'd23;    
		mem[  1666] = 10'd37;    
		mem[  1667] = 10'd27;    
		mem[  1668] = 10'd30;    
		mem[  1669] = 10'd66;    
		mem[  1670] = 10'd26;    
		mem[  1671] = 10'd65;    
		mem[  1672] = 10'd31;    
		mem[  1673] = 10'd60;    
		mem[  1674] = 10'd31;    
		mem[  1675] = 10'd22;    
		mem[  1676] = 10'd41;    
		mem[  1677] = 10'd24;    
		mem[  1678] = 10'd30;    
		mem[  1679] = 10'd32;    
		mem[  1680] = 10'd36;    
		mem[  1681] = 10'd25;    
		mem[  1682] = 10'd33;    
		mem[  1683] = 10'd32;    
		mem[  1684] = 10'd29;    
		mem[  1685] = 10'd65;    
		mem[  1686] = 10'd28;    
		mem[  1687] = 10'd64;    
		mem[  1688] = 10'd21;    
		mem[  1689] = 10'd33;    
		mem[  1690] = 10'd35;    
		mem[  1691] = 10'd33;    
		mem[  1692] = 10'd25;    
		mem[  1693] = 10'd36;    
		mem[  1694] = 10'd28;    
		mem[  1695] = 10'd29;    
		mem[  1696] = 10'd30;    
		mem[  1697] = 10'd37;    
		mem[  1698] = 10'd26;    
		mem[  1699] = 10'd29;    
		mem[  1700] = 10'd35;    
		mem[  1701] = 10'd31;    
		mem[  1702] = 10'd25;    
		mem[  1703] = 10'd33;    
		mem[  1704] = 10'd30;    
		mem[  1705] = 10'd24;    
		mem[  1706] = 10'd34;    
		mem[  1707] = 10'd27;    
		mem[  1708] = 10'd28;    
		mem[  1709] = 10'd27;    
		mem[  1710] = 10'd35;    
		mem[  1711] = 10'd27;    
		mem[  1712] = 10'd24;    
		mem[  1713] = 10'd36;    
		mem[  1714] = 10'd24;    
		mem[  1715] = 10'd29;    
		mem[  1716] = 10'd29;    
		mem[  1717] = 10'd33;    
		mem[  1718] = 10'd26;    
		mem[  1719] = 10'd27;    
		mem[  1720] = 10'd34;    
		mem[  1721] = 10'd26;    
		mem[  1722] = 10'd27;    
		mem[  1723] = 10'd31;    
		mem[  1724] = 10'd32;    
		mem[  1725] = 10'd25;    
		mem[  1726] = 10'd30;    
		mem[  1727] = 10'd31;    
		mem[  1728] = 10'd29;    
		mem[  1729] = 10'd25;    
		mem[  1730] = 10'd33;    
		mem[  1731] = 10'd29;    
		mem[  1732] = 10'd25;    
		mem[  1733] = 10'd33;    
		mem[  1734] = 10'd27;    
		mem[  1735] = 10'd29;    
		mem[  1736] = 10'd27;    
		mem[  1737] = 10'd34;    
		mem[  1738] = 10'd27;    
		mem[  1739] = 10'd25;    
		mem[  1740] = 10'd34;    
		mem[  1741] = 10'd26;    
		mem[  1742] = 10'd29;    
		mem[  1743] = 10'd29;    
		mem[  1744] = 10'd32;    
		mem[  1745] = 10'd27;    
		mem[  1746] = 10'd28;    
		mem[  1747] = 10'd32;    
		mem[  1748] = 10'd27;    
		mem[  1749] = 10'd28;    
		mem[  1750] = 10'd30;    
		mem[  1751] = 10'd31;    
		mem[  1752] = 10'd26;    
		mem[  1753] = 10'd28;    
		mem[  1754] = 10'd29;    
		mem[  1755] = 10'd26;    
		mem[  1756] = 10'd26;    
		mem[  1757] = 10'd28;    
		mem[  1758] = 10'd29;    
		mem[  1759] = 10'd26;    
		mem[  1760] = 10'd27;    
		mem[  1761] = 10'd29;    
		mem[  1762] = 10'd25;    
		mem[  1763] = 10'd27;    
		mem[  1764] = 10'd28;    
		mem[  1765] = 10'd30;    
		mem[  1766] = 10'd25;    
		mem[  1767] = 10'd26;    
		mem[  1768] = 10'd30;    
		mem[  1769] = 10'd25;    
		mem[  1770] = 10'd28;    
		mem[  1771] = 10'd27;    
		mem[  1772] = 10'd29;    
		mem[  1773] = 10'd27;    
		mem[  1774] = 10'd25;    
		mem[  1775] = 10'd30;    
		mem[  1776] = 10'd26;    
		mem[  1777] = 10'd27;    
		mem[  1778] = 10'd27;    
		mem[  1779] = 10'd29;    
		mem[  1780] = 10'd27;    
		mem[  1781] = 10'd26;    
		mem[  1782] = 10'd29;    
		mem[  1783] = 10'd27;    
		mem[  1784] = 10'd27;    
		mem[  1785] = 10'd26;    
		mem[  1786] = 10'd29;    
		mem[  1787] = 10'd28;    
		mem[  1788] = 10'd25;    
		mem[  1789] = 10'd29;    
		mem[  1790] = 10'd27;    
		mem[  1791] = 10'd28;    
		mem[  1792] = 10'd25;    
		mem[  1793] = 10'd29;    
		mem[  1794] = 10'd28;    
		mem[  1795] = 10'd26;    
		mem[  1796] = 10'd27;    
		mem[  1797] = 10'd28;    
		mem[  1798] = 10'd27;    
		mem[  1799] = 10'd27;    
		mem[  1800] = 10'd28;    
		mem[  1801] = 10'd28;    
		mem[  1802] = 10'd26;    
		mem[  1803] = 10'd27;    
		mem[  1804] = 10'd29;    
		mem[  1805] = 10'd26;    
		mem[  1806] = 10'd213;    
		mem[  1807] = 10'd106;    
		mem[  1808] = 10'd68;    
		mem[  1809] = 10'd132;    
		mem[  1810] = 10'd192;    
		mem[  1811] = 10'd776;    
		mem[  1812] = 10'd57;    
		mem[  1813] = 10'd24;    
		mem[  1814] = 10'd23;    
		mem[  1815] = 10'd35;    
		mem[  1816] = 10'd23;    
		mem[  1817] = 10'd58;    
		mem[  1818] = 10'd18;    
		mem[  1819] = 10'd28;    
		mem[  1820] = 10'd32;    
		mem[  1821] = 10'd30;    
		mem[  1822] = 10'd21;    
		mem[  1823] = 10'd32;    
		mem[  1824] = 10'd25;    
		mem[  1825] = 10'd27;    
		mem[  1826] = 10'd59;    
		mem[  1827] = 10'd24;    
		mem[  1828] = 10'd57;    
		mem[  1829] = 10'd28;    
		mem[  1830] = 10'd20;    
		mem[  1831] = 10'd33;    
		mem[  1832] = 10'd28;    
		mem[  1833] = 10'd20;    
		mem[  1834] = 10'd36;    
		mem[  1835] = 10'd22;    
		mem[  1836] = 10'd27;    
		mem[  1837] = 10'd28;    
		mem[  1838] = 10'd32;    
		mem[  1839] = 10'd22;    
		mem[  1840] = 10'd30;    
		mem[  1841] = 10'd28;    
		mem[  1842] = 10'd26;    
		mem[  1843] = 10'd23;    
		mem[  1844] = 10'd35;    
		mem[  1845] = 10'd25;    
		mem[  1846] = 10'd56;    
		mem[  1847] = 10'd25;    
		mem[  1848] = 10'd24;    
		mem[  1849] = 10'd31;    
		mem[  1850] = 10'd29;    
		mem[  1851] = 10'd22;    
		mem[  1852] = 10'd33;    
		mem[  1853] = 10'd24;    
		mem[  1854] = 10'd27;    
		mem[  1855] = 10'd27;    
		mem[  1856] = 10'd32;    
		mem[  1857] = 10'd24;    
		mem[  1858] = 10'd26;    
		mem[  1859] = 10'd30;    
		mem[  1860] = 10'd26;    
		mem[  1861] = 10'd21;    
		mem[  1862] = 10'd30;    
		mem[  1863] = 10'd27;    
		mem[  1864] = 10'd21;    
		mem[  1865] = 10'd30;    
		mem[  1866] = 10'd24;    
		mem[  1867] = 10'd26;    
		mem[  1868] = 10'd23;    
		mem[  1869] = 10'd31;    
		mem[  1870] = 10'd24;    
		mem[  1871] = 10'd22;    
		mem[  1872] = 10'd32;    
		mem[  1873] = 10'd22;    
		mem[  1874] = 10'd25;    
		mem[  1875] = 10'd26;    
		mem[  1876] = 10'd30;    
		mem[  1877] = 10'd23;    
		mem[  1878] = 10'd23;    
		mem[  1879] = 10'd31;    
		mem[  1880] = 10'd20;    
		mem[  1881] = 10'd27;    
		mem[  1882] = 10'd27;    
		mem[  1883] = 10'd29;    
		mem[  1884] = 10'd23;    
		mem[  1885] = 10'd25;    
		mem[  1886] = 10'd29;    
		mem[  1887] = 10'd26;    
		mem[  1888] = 10'd22;    
		mem[  1889] = 10'd29;    
		mem[  1890] = 10'd26;    
		mem[  1891] = 10'd22;    
		mem[  1892] = 10'd29;    
		mem[  1893] = 10'd25;    
		mem[  1894] = 10'd26;    
		mem[  1895] = 10'd23;    
		mem[  1896] = 10'd30;    
		mem[  1897] = 10'd25;    
		mem[  1898] = 10'd22;    
		mem[  1899] = 10'd31;    
		mem[  1900] = 10'd23;    
		mem[  1901] = 10'd25;    
		mem[  1902] = 10'd26;    
		mem[  1903] = 10'd28;    
		mem[  1904] = 10'd25;    
		mem[  1905] = 10'd24;    
		mem[  1906] = 10'd29;    
		mem[  1907] = 10'd24;    
		mem[  1908] = 10'd25;    
		mem[  1909] = 10'd26;    
		mem[  1910] = 10'd28;    
		mem[  1911] = 10'd24;    
		mem[  1912] = 10'd26;    
		mem[  1913] = 10'd27;    
		mem[  1914] = 10'd26;    
		mem[  1915] = 10'd23;    
		mem[  1916] = 10'd27;    
		mem[  1917] = 10'd25;    
		mem[  1918] = 10'd22;    
		mem[  1919] = 10'd26;    
		mem[  1920] = 10'd25;    
		mem[  1921] = 10'd25;    
		mem[  1922] = 10'd22;    
		mem[  1923] = 10'd26;    
		mem[  1924] = 10'd26;    
		mem[  1925] = 10'd22;    
		mem[  1926] = 10'd24;    
		mem[  1927] = 10'd27;    
		mem[  1928] = 10'd23;    
		mem[  1929] = 10'd23;    
		mem[  1930] = 10'd26;    
		mem[  1931] = 10'd26;    
		mem[  1932] = 10'd23;    
		mem[  1933] = 10'd24;    
		mem[  1934] = 10'd26;    
		mem[  1935] = 10'd23;    
		mem[  1936] = 10'd24;    
		mem[  1937] = 10'd25;    
		mem[  1938] = 10'd26;    
		mem[  1939] = 10'd23;    
		mem[  1940] = 10'd24;    
		mem[  1941] = 10'd26;    
		mem[  1942] = 10'd22;    
		mem[  1943] = 10'd25;    
		mem[  1944] = 10'd25;    
		mem[  1945] = 10'd26;    
		mem[  1946] = 10'd24;    
		mem[  1947] = 10'd23;    
		mem[  1948] = 10'd26;    
		mem[  1949] = 10'd23;    
		mem[  1950] = 10'd25;    
		mem[  1951] = 10'd24;    
		mem[  1952] = 10'd26;    
		mem[  1953] = 10'd24;    
		mem[  1954] = 10'd23;    
		mem[  1955] = 10'd26;    
		mem[  1956] = 10'd24;    
		mem[  1957] = 10'd24;    
		mem[  1958] = 10'd24;    
		mem[  1959] = 10'd26;    
		mem[  1960] = 10'd24;    
		mem[  1961] = 10'd24;    
		mem[  1962] = 10'd25;    
		mem[  1963] = 10'd25;    
		mem[  1964] = 10'd24;    
		mem[  1965] = 10'd24;    
		mem[  1966] = 10'd25;    
		mem[  1967] = 10'd25;    
		mem[  1968] = 10'd23;    
		mem[  1969] = 10'd25;    
		mem[  1970] = 10'd25;    
		mem[  1971] = 10'd25;    
		mem[  1972] = 10'd23;    
		mem[  1973] = 10'd25;    
		mem[  1974] = 10'd25;    
		mem[  1975] = 10'd193;    
		mem[  1976] = 10'd1023;// 10'd1305;    
		mem[  1977] = 10'd44;    
		mem[  1978] = 10'd22;    
		mem[  1979] = 10'd17;    
		mem[  1980] = 10'd45;    
		mem[  1981] = 10'd16;    
		mem[  1982] = 10'd21;    
		mem[  1983] = 10'd44;    
		mem[  1984] = 10'd22;    
		mem[  1985] = 10'd16;    
		mem[  1986] = 10'd20;    
		mem[  1987] = 10'd26;    
		mem[  1988] = 10'd15;    
		mem[  1989] = 10'd21;    
		mem[  1990] = 10'd19;    
		mem[  1991] = 10'd25;    
		mem[  1992] = 10'd22;    
		mem[  1993] = 10'd16;    
		mem[  1994] = 10'd20;    
		mem[  1995] = 10'd26;    
		mem[  1996] = 10'd15;    
		mem[  1997] = 10'd21;    
		mem[  1998] = 10'd19;    
		mem[  1999] = 10'd25;    
		mem[  2000] = 10'd21;    
		mem[  2001] = 10'd17;    
		mem[  2002] = 10'd20;    
		mem[  2003] = 10'd25;    
		mem[  2004] = 10'd16;    
		mem[  2005] = 10'd21;    
		mem[  2006] = 10'd18;    
		mem[  2007] = 10'd26;    
		mem[  2008] = 10'd21;    
		mem[  2009] = 10'd17;    
		mem[  2010] = 10'd19;    
		mem[  2011] = 10'd26;    
		mem[  2012] = 10'd16;    
		mem[  2013] = 10'd21;    
		mem[  2014] = 10'd18;    
		mem[  2015] = 10'd25;    
		mem[  2016] = 10'd22;    
		mem[  2017] = 10'd16;    
		mem[  2018] = 10'd20;    
		mem[  2019] = 10'd25;    
		mem[  2020] = 10'd16;    
		mem[  2021] = 10'd21;    
		mem[  2022] = 10'd19;    
		mem[  2023] = 10'd25;    
		mem[  2024] = 10'd21;    
		mem[  2025] = 10'd17;    
		mem[  2026] = 10'd20;    
		mem[  2027] = 10'd25;    
		mem[  2028] = 10'd16;    
		mem[  2029] = 10'd21;    
		mem[  2030] = 10'd19;    
		mem[  2031] = 10'd25;    
		mem[  2032] = 10'd21;    
		mem[  2033] = 10'd17;    
		mem[  2034] = 10'd20;    
		mem[  2035] = 10'd25;    
		mem[  2036] = 10'd16;    
		mem[  2037] = 10'd21;    
		mem[  2038] = 10'd19;    
		mem[  2039] = 10'd24;    
		mem[  2040] = 10'd22;    
		mem[  2041] = 10'd17;    
		mem[  2042] = 10'd20;    
		mem[  2043] = 10'd24;    
		mem[  2044] = 10'd17;    
		mem[  2045] = 10'd21;    
		mem[  2046] = 10'd19;    
		mem[  2047] = 10'd24;    
		mem[  2048] = 10'd21;    
		mem[  2049] = 10'd18;    
		mem[  2050] = 10'd20;    
		mem[  2051] = 10'd24;    
		mem[  2052] = 10'd17;    
		mem[  2053] = 10'd21;    
		mem[  2054] = 10'd19;    
		mem[  2055] = 10'd24;    
		mem[  2056] = 10'd21;    
		mem[  2057] = 10'd18;    
		mem[  2058] = 10'd20;    
		mem[  2059] = 10'd24;    
		mem[  2060] = 10'd17;    
		mem[  2061] = 10'd21;    
		mem[  2062] = 10'd19;    
		mem[  2063] = 10'd24;    
		mem[  2064] = 10'd21;    
		mem[  2065] = 10'd17;    
		mem[  2066] = 10'd21;    
		mem[  2067] = 10'd24;    
		mem[  2068] = 10'd17;    
		mem[  2069] = 10'd21;    
		mem[  2070] = 10'd19;    
		mem[  2071] = 10'd23;    
		mem[  2072] = 10'd22;    
		mem[  2073] = 10'd17;    
		mem[  2074] = 10'd20;    
		mem[  2075] = 10'd24;    
		mem[  2076] = 10'd17;    
		mem[  2077] = 10'd21;    
		mem[  2078] = 10'd20;    
		mem[  2079] = 10'd23;    
		mem[  2080] = 10'd21;    
		mem[  2081] = 10'd18;    
		mem[  2082] = 10'd21;    
		mem[  2083] = 10'd23;    
		mem[  2084] = 10'd17;    
		mem[  2085] = 10'd21;    
		mem[  2086] = 10'd20;    
		mem[  2087] = 10'd23;    
		mem[  2088] = 10'd21;    
		mem[  2089] = 10'd18;    
		mem[  2090] = 10'd20;    
		mem[  2091] = 10'd24;    
		mem[  2092] = 10'd17;    
		mem[  2093] = 10'd21;    
		mem[  2094] = 10'd20;    
		mem[  2095] = 10'd23;    
		mem[  2096] = 10'd21;    
		mem[  2097] = 10'd18;    
		mem[  2098] = 10'd20;    
		mem[  2099] = 10'd23;    
		mem[  2100] = 10'd18;    
		mem[  2101] = 10'd21;    
		mem[  2102] = 10'd20;    
		mem[  2103] = 10'd23;    
		mem[  2104] = 10'd20;    
		mem[  2105] = 10'd19;    
		mem[  2106] = 10'd20;    
		mem[  2107] = 10'd23;    
		mem[  2108] = 10'd18;    
		mem[  2109] = 10'd21;    
		mem[  2110] = 10'd20;    
		mem[  2111] = 10'd22;    
		mem[  2112] = 10'd21;    
		mem[  2113] = 10'd19;    
		mem[  2114] = 10'd20;    
		mem[  2115] = 10'd138;    
		mem[  2116] = 10'd65;    
		mem[  2117] = 10'd20;    
		mem[  2118] = 10'd83;    
		mem[  2119] = 10'd61;    
		mem[  2120] = 10'd22;    
		mem[  2121] = 10'd80;    
		mem[  2122] = 10'd62;    
		mem[  2123] = 10'd21;    
		mem[  2124] = 10'd81;    
		mem[  2125] = 10'd62;    
		mem[  2126] = 10'd22;    
		mem[  2127] = 10'd78;    
		mem[  2128] = 10'd63;    
		mem[  2129] = 10'd21;    
		mem[  2130] = 10'd82;    
		mem[  2131] = 10'd61;    
		mem[  2132] = 10'd21;    
		mem[  2133] = 10'd79;    
		mem[  2134] = 10'd63;    
		mem[  2135] = 10'd21;    
		mem[  2136] = 10'd83;    
		mem[  2137] = 10'd60;    
		mem[  2138] = 10'd22;    
		mem[  2139] = 10'd80;    
		mem[  2140] = 10'd60;    
		mem[  2141] = 10'd20;    
		mem[  2142] = 10'd86;    
		mem[  2143] = 10'd61;    
		mem[  2144] = 10'd21;    
		mem[  2145] = 10'd80;    
		mem[  2146] = 10'd58;    
		mem[  2147] = 10'd170;    
		mem[  2148] = 10'd20;    
		mem[  2149] = 10'd78;    
		mem[  2150] = 10'd64;    
		mem[  2151] = 10'd19;    
		mem[  2152] = 10'd1023;    
		mem[  2153] = 10'd1023;    
	end
	
endmodule

