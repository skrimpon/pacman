module pacman_wakka(in, out, clk);
	 input [11:0] in;
	 input clk;
	 output reg [10:0] out;
	 
	 reg  [10:0] mem [0:2834];
	 always @(posedge clk) out  =  mem[ in ];
	 
	 initial begin
		mem[     0] = 11'd2001;    
		mem[     1] = 11'd31;    
		mem[     2] = 11'd61;    
		mem[     3] = 11'd22;    
		mem[     4] = 11'd113;    
		mem[     5] = 11'd65;    
		mem[     6] = 11'd33;    
		mem[     7] = 11'd33;    
		mem[     8] = 11'd63;    
		mem[     9] = 11'd64;    
		mem[    10] = 11'd68;    
		mem[    11] = 11'd28;    
		mem[    12] = 11'd33;    
		mem[    13] = 11'd68;    
		mem[    14] = 11'd31;    
		mem[    15] = 11'd26;    
		mem[    16] = 11'd65;    
		mem[    17] = 11'd58;    
		mem[    18] = 11'd65;    
		mem[    19] = 11'd58;    
		mem[    20] = 11'd64;    
		mem[    21] = 11'd58;    
		mem[    22] = 11'd65;    
		mem[    23] = 11'd58;    
		mem[    24] = 11'd64;    
		mem[    25] = 11'd59;    
		mem[    26] = 11'd64;    
		mem[    27] = 11'd32;    
		mem[    28] = 11'd26;    
		mem[    29] = 11'd64;    
		mem[    30] = 11'd59;    
		mem[    31] = 11'd64;    
		mem[    32] = 11'd32;    
		mem[    33] = 11'd26;    
		mem[    34] = 11'd64;    
		mem[    35] = 11'd59;    
		mem[    36] = 11'd64;    
		mem[    37] = 11'd32;    
		mem[    38] = 11'd26;    
		mem[    39] = 11'd31;    
		mem[    40] = 11'd33;    
		mem[    41] = 11'd59;    
		mem[    42] = 11'd64;    
		mem[    43] = 11'd32;    
		mem[    44] = 11'd27;    
		mem[    45] = 11'd30;    
		mem[    46] = 11'd33;    
		mem[    47] = 11'd59;    
		mem[    48] = 11'd64;    
		mem[    49] = 11'd32;    
		mem[    50] = 11'd27;    
		mem[    51] = 11'd31;    
		mem[    52] = 11'd32;    
		mem[    53] = 11'd60;    
		mem[    54] = 11'd63;    
		mem[    55] = 11'd32;    
		mem[    56] = 11'd27;    
		mem[    57] = 11'd31;    
		mem[    58] = 11'd32;    
		mem[    59] = 11'd60;    
		mem[    60] = 11'd60;    
		mem[    61] = 11'd62;    
		mem[    62] = 11'd31;    
		mem[    63] = 11'd31;    
		mem[    64] = 11'd32;    
		mem[    65] = 11'd30;    
		mem[    66] = 11'd31;    
		mem[    67] = 11'd30;    
		mem[    68] = 11'd31;    
		mem[    69] = 11'd30;    
		mem[    70] = 11'd32;    
		mem[    71] = 11'd30;    
		mem[    72] = 11'd31;    
		mem[    73] = 11'd30;    
		mem[    74] = 11'd31;    
		mem[    75] = 11'd30;    
		mem[    76] = 11'd31;    
		mem[    77] = 11'd30;    
		mem[    78] = 11'd32;    
		mem[    79] = 11'd29;    
		mem[    80] = 11'd32;    
		mem[    81] = 11'd30;    
		mem[    82] = 11'd32;    
		mem[    83] = 11'd32;    
		mem[    84] = 11'd33;    
		mem[    85] = 11'd31;    
		mem[    86] = 11'd34;    
		mem[    87] = 11'd32;    
		mem[    88] = 11'd33;    
		mem[    89] = 11'd31;    
		mem[    90] = 11'd33;    
		mem[    91] = 11'd32;    
		mem[    92] = 11'd34;    
		mem[    93] = 11'd32;    
		mem[    94] = 11'd33;    
		mem[    95] = 11'd31;    
		mem[    96] = 11'd33;    
		mem[    97] = 11'd32;    
		mem[    98] = 11'd34;    
		mem[    99] = 11'd31;    
		mem[   100] = 11'd34;    
		mem[   101] = 11'd31;    
		mem[   102] = 11'd33;    
		mem[   103] = 11'd32;    
		mem[   104] = 11'd33;    
		mem[   105] = 11'd30;    
		mem[   106] = 11'd31;    
		mem[   107] = 11'd30;    
		mem[   108] = 11'd31;    
		mem[   109] = 11'd31;    
		mem[   110] = 11'd31;    
		mem[   111] = 11'd30;    
		mem[   112] = 11'd31;    
		mem[   113] = 11'd30;    
		mem[   114] = 11'd31;    
		mem[   115] = 11'd31;    
		mem[   116] = 11'd31;    
		mem[   117] = 11'd30;    
		mem[   118] = 11'd31;    
		mem[   119] = 11'd30;    
		mem[   120] = 11'd31;    
		mem[   121] = 11'd30;    
		mem[   122] = 11'd32;    
		mem[   123] = 11'd30;    
		mem[   124] = 11'd31;    
		mem[   125] = 11'd30;    
		mem[   126] = 11'd31;    
		mem[   127] = 11'd30;    
		mem[   128] = 11'd32;    
		mem[   129] = 11'd89;    
		mem[   130] = 11'd65;    
		mem[   131] = 11'd58;    
		mem[   132] = 11'd64;    
		mem[   133] = 11'd32;    
		mem[   134] = 11'd25;    
		mem[   135] = 11'd66;    
		mem[   136] = 11'd58;    
		mem[   137] = 11'd64;    
		mem[   138] = 11'd58;    
		mem[   139] = 11'd65;    
		mem[   140] = 11'd58;    
		mem[   141] = 11'd64;    
		mem[   142] = 11'd33;    
		mem[   143] = 11'd25;    
		mem[   144] = 11'd65;    
		mem[   145] = 11'd58;    
		mem[   146] = 11'd65;    
		mem[   147] = 11'd57;    
		mem[   148] = 11'd65;    
		mem[   149] = 11'd58;    
		mem[   150] = 11'd64;    
		mem[   151] = 11'd59;    
		mem[   152] = 11'd64;    
		mem[   153] = 11'd58;    
		mem[   154] = 11'd62;    
		mem[   155] = 11'd30;    
		mem[   156] = 11'd32;    
		mem[   157] = 11'd30;    
		mem[   158] = 11'd31;    
		mem[   159] = 11'd32;    
		mem[   160] = 11'd30;    
		mem[   161] = 11'd31;    
		mem[   162] = 11'd30;    
		mem[   163] = 11'd32;    
		mem[   164] = 11'd30;    
		mem[   165] = 11'd31;    
		mem[   166] = 11'd30;    
		mem[   167] = 11'd31;    
		mem[   168] = 11'd30;    
		mem[   169] = 11'd31;    
		mem[   170] = 11'd30;    
		mem[   171] = 11'd32;    
		mem[   172] = 11'd30;    
		mem[   173] = 11'd31;    
		mem[   174] = 11'd30;    
		mem[   175] = 11'd31;    
		mem[   176] = 11'd30;    
		mem[   177] = 11'd36;    
		mem[   178] = 11'd64;    
		mem[   179] = 11'd15;    
		mem[   180] = 11'd79;    
		mem[   181] = 11'd33;    
		mem[   182] = 11'd99;    
		mem[   183] = 11'd28;    
		mem[   184] = 11'd34;    
		mem[   185] = 11'd58;    
		mem[   186] = 11'd22;    
		mem[   187] = 11'd50;    
		mem[   188] = 11'd67;    
		mem[   189] = 11'd66;    
		mem[   190] = 11'd32;    
		mem[   191] = 11'd32;    
		mem[   192] = 11'd62;    
		mem[   193] = 11'd61;    
		mem[   194] = 11'd63;    
		mem[   195] = 11'd29;    
		mem[   196] = 11'd30;    
		mem[   197] = 11'd62;    
		mem[   198] = 11'd61;    
		mem[   199] = 11'd63;    
		mem[   200] = 11'd29;    
		mem[   201] = 11'd30;    
		mem[   202] = 11'd62;    
		mem[   203] = 11'd61;    
		mem[   204] = 11'd63;    
		mem[   205] = 11'd29;    
		mem[   206] = 11'd31;    
		mem[   207] = 11'd61;    
		mem[   208] = 11'd61;    
		mem[   209] = 11'd63;    
		mem[   210] = 11'd14;    
		mem[   211] = 11'd15;    
		mem[   212] = 11'd31;    
		mem[   213] = 11'd61;    
		mem[   214] = 11'd61;    
		mem[   215] = 11'd63;    
		mem[   216] = 11'd14;    
		mem[   217] = 11'd15;    
		mem[   218] = 11'd31;    
		mem[   219] = 11'd61;    
		mem[   220] = 11'd61;    
		mem[   221] = 11'd63;    
		mem[   222] = 11'd14;    
		mem[   223] = 11'd15;    
		mem[   224] = 11'd31;    
		mem[   225] = 11'd61;    
		mem[   226] = 11'd61;    
		mem[   227] = 11'd63;    
		mem[   228] = 11'd29;    
		mem[   229] = 11'd31;    
		mem[   230] = 11'd62;    
		mem[   231] = 11'd60;    
		mem[   232] = 11'd63;    
		mem[   233] = 11'd30;    
		mem[   234] = 11'd30;    
		mem[   235] = 11'd62;    
		mem[   236] = 11'd61;    
		mem[   237] = 11'd62;    
		mem[   238] = 11'd30;    
		mem[   239] = 11'd33;    
		mem[   240] = 11'd59;    
		mem[   241] = 11'd32;    
		mem[   242] = 11'd29;    
		mem[   243] = 11'd31;    
		mem[   244] = 11'd30;    
		mem[   245] = 11'd30;    
		mem[   246] = 11'd31;    
		mem[   247] = 11'd30;    
		mem[   248] = 11'd31;    
		mem[   249] = 11'd30;    
		mem[   250] = 11'd31;    
		mem[   251] = 11'd30;    
		mem[   252] = 11'd31;    
		mem[   253] = 11'd31;    
		mem[   254] = 11'd31;    
		mem[   255] = 11'd30;    
		mem[   256] = 11'd31;    
		mem[   257] = 11'd31;    
		mem[   258] = 11'd30;    
		mem[   259] = 11'd31;    
		mem[   260] = 11'd31;    
		mem[   261] = 11'd30;    
		mem[   262] = 11'd33;    
		mem[   263] = 11'd40;    
		mem[   264] = 11'd38;    
		mem[   265] = 11'd40;    
		mem[   266] = 11'd38;    
		mem[   267] = 11'd39;    
		mem[   268] = 11'd39;    
		mem[   269] = 11'd39;    
		mem[   270] = 11'd38;    
		mem[   271] = 11'd40;    
		mem[   272] = 11'd38;    
		mem[   273] = 11'd40;    
		mem[   274] = 11'd38;    
		mem[   275] = 11'd39;    
		mem[   276] = 11'd39;    
		mem[   277] = 11'd39;    
		mem[   278] = 11'd38;    
		mem[   279] = 11'd40;    
		mem[   280] = 11'd38;    
		mem[   281] = 11'd40;    
		mem[   282] = 11'd35;    
		mem[   283] = 11'd37;    
		mem[   284] = 11'd35;    
		mem[   285] = 11'd37;    
		mem[   286] = 11'd36;    
		mem[   287] = 11'd38;    
		mem[   288] = 11'd36;    
		mem[   289] = 11'd37;    
		mem[   290] = 11'd36;    
		mem[   291] = 11'd36;    
		mem[   292] = 11'd37;    
		mem[   293] = 11'd37;    
		mem[   294] = 11'd36;    
		mem[   295] = 11'd37;    
		mem[   296] = 11'd36;    
		mem[   297] = 11'd38;    
		mem[   298] = 11'd36;    
		mem[   299] = 11'd37;    
		mem[   300] = 11'd36;    
		mem[   301] = 11'd144;    
		mem[   302] = 11'd77;    
		mem[   303] = 11'd39;    
		mem[   304] = 11'd30;    
		mem[   305] = 11'd78;    
		mem[   306] = 11'd73;    
		mem[   307] = 11'd35;    
		mem[   308] = 11'd36;    
		mem[   309] = 11'd76;    
		mem[   310] = 11'd36;    
		mem[   311] = 11'd17;    
		mem[   312] = 11'd87;    
		mem[   313] = 11'd21;    
		mem[   314] = 11'd64;    
		mem[   315] = 11'd77;    
		mem[   316] = 11'd83;    
		mem[   317] = 11'd21;    
		mem[   318] = 11'd65;    
		mem[   319] = 11'd78;    
		mem[   320] = 11'd81;    
		mem[   321] = 11'd21;    
		mem[   322] = 11'd65;    
		mem[   323] = 11'd46;    
		mem[   324] = 11'd21;    
		mem[   325] = 11'd12;    
		mem[   326] = 11'd81;    
		mem[   327] = 11'd84;    
		mem[   328] = 11'd41;    
		mem[   329] = 11'd42;    
		mem[   330] = 11'd42;    
		mem[   331] = 11'd40;    
		mem[   332] = 11'd43;    
		mem[   333] = 11'd39;    
		mem[   334] = 11'd43;    
		mem[   335] = 11'd39;    
		mem[   336] = 11'd43;    
		mem[   337] = 11'd39;    
		mem[   338] = 11'd42;    
		mem[   339] = 11'd40;    
		mem[   340] = 11'd42;    
		mem[   341] = 11'd40;    
		mem[   342] = 11'd42;    
		mem[   343] = 11'd57;    
		mem[   344] = 11'd12;    
		mem[   345] = 11'd30;    
		mem[   346] = 11'd63;    
		mem[   347] = 11'd60;    
		mem[   348] = 11'd34;    
		mem[   349] = 11'd14;    
		mem[   350] = 11'd13;    
		mem[   351] = 11'd60;    
		mem[   352] = 11'd64;    
		mem[   353] = 11'd60;    
		mem[   354] = 11'd34;    
		mem[   355] = 11'd14;    
		mem[   356] = 11'd13;    
		mem[   357] = 11'd60;    
		mem[   358] = 11'd64;    
		mem[   359] = 11'd60;    
		mem[   360] = 11'd34;    
		mem[   361] = 11'd14;    
		mem[   362] = 11'd13;    
		mem[   363] = 11'd60;    
		mem[   364] = 11'd64;    
		mem[   365] = 11'd60;    
		mem[   366] = 11'd34;    
		mem[   367] = 11'd14;    
		mem[   368] = 11'd13;    
		mem[   369] = 11'd60;    
		mem[   370] = 11'd64;    
		mem[   371] = 11'd60;    
		mem[   372] = 11'd34;    
		mem[   373] = 11'd14;    
		mem[   374] = 11'd13;    
		mem[   375] = 11'd60;    
		mem[   376] = 11'd63;    
		mem[   377] = 11'd61;    
		mem[   378] = 11'd34;    
		mem[   379] = 11'd14;    
		mem[   380] = 11'd32;    
		mem[   381] = 11'd115;    
		mem[   382] = 11'd91;    
		mem[   383] = 11'd32;    
		mem[   384] = 11'd121;    
		mem[   385] = 11'd92;    
		mem[   386] = 11'd32;    
		mem[   387] = 11'd121;    
		mem[   388] = 11'd93;    
		mem[   389] = 11'd7;    
		mem[   390] = 11'd65;    
		mem[   391] = 11'd35;    
		mem[   392] = 11'd29;    
		mem[   393] = 11'd60;    
		mem[   394] = 11'd35;    
		mem[   395] = 11'd25;    
		mem[   396] = 11'd31;    
		mem[   397] = 11'd31;    
		mem[   398] = 11'd63;    
		mem[   399] = 11'd28;    
		mem[   400] = 11'd32;    
		mem[   401] = 11'd35;    
		mem[   402] = 11'd25;    
		mem[   403] = 11'd32;    
		mem[   404] = 11'd18;    
		mem[   405] = 11'd12;    
		mem[   406] = 11'd35;    
		mem[   407] = 11'd28;    
		mem[   408] = 11'd29;    
		mem[   409] = 11'd31;    
		mem[   410] = 11'd34;    
		mem[   411] = 11'd30;    
		mem[   412] = 11'd60;    
		mem[   413] = 11'd31;    
		mem[   414] = 11'd30;    
		mem[   415] = 11'd31;    
		mem[   416] = 11'd29;    
		mem[   417] = 11'd31;    
		mem[   418] = 11'd31;    
		mem[   419] = 11'd30;    
		mem[   420] = 11'd31;    
		mem[   421] = 11'd30;    
		mem[   422] = 11'd31;    
		mem[   423] = 11'd30;    
		mem[   424] = 11'd31;    
		mem[   425] = 11'd31;    
		mem[   426] = 11'd31;    
		mem[   427] = 11'd30;    
		mem[   428] = 11'd31;    
		mem[   429] = 11'd31;    
		mem[   430] = 11'd30;    
		mem[   431] = 11'd31;    
		mem[   432] = 11'd31;    
		mem[   433] = 11'd30;    
		mem[   434] = 11'd31;    
		mem[   435] = 11'd31;    
		mem[   436] = 11'd30;    
		mem[   437] = 11'd31;    
		mem[   438] = 11'd31;    
		mem[   439] = 11'd31;    
		mem[   440] = 11'd30;    
		mem[   441] = 11'd31;    
		mem[   442] = 11'd30;    
		mem[   443] = 11'd31;    
		mem[   444] = 11'd30;    
		mem[   445] = 11'd31;    
		mem[   446] = 11'd30;    
		mem[   447] = 11'd31;    
		mem[   448] = 11'd31;    
		mem[   449] = 11'd31;    
		mem[   450] = 11'd30;    
		mem[   451] = 11'd31;    
		mem[   452] = 11'd30;    
		mem[   453] = 11'd31;    
		mem[   454] = 11'd31;    
		mem[   455] = 11'd31;    
		mem[   456] = 11'd30;    
		mem[   457] = 11'd32;    
		mem[   458] = 11'd30;    
		mem[   459] = 11'd31;    
		mem[   460] = 11'd30;    
		mem[   461] = 11'd31;    
		mem[   462] = 11'd30;    
		mem[   463] = 11'd31;    
		mem[   464] = 11'd30;    
		mem[   465] = 11'd31;    
		mem[   466] = 11'd30;    
		mem[   467] = 11'd31;    
		mem[   468] = 11'd31;    
		mem[   469] = 11'd30;    
		mem[   470] = 11'd31;    
		mem[   471] = 11'd31;    
		mem[   472] = 11'd30;    
		mem[   473] = 11'd31;    
		mem[   474] = 11'd30;    
		mem[   475] = 11'd31;    
		mem[   476] = 11'd31;    
		mem[   477] = 11'd30;    
		mem[   478] = 11'd31;    
		mem[   479] = 11'd31;    
		mem[   480] = 11'd30;    
		mem[   481] = 11'd27;    
		mem[   482] = 11'd28;    
		mem[   483] = 11'd105;    
		mem[   484] = 11'd23;    
		mem[   485] = 11'd80;    
		mem[   486] = 11'd49;    
		mem[   487] = 11'd52;    
		mem[   488] = 11'd53;    
		mem[   489] = 11'd50;    
		mem[   490] = 11'd52;    
		mem[   491] = 11'd30;    
		mem[   492] = 11'd20;    
		mem[   493] = 11'd55;    
		mem[   494] = 11'd50;    
		mem[   495] = 11'd53;    
		mem[   496] = 11'd46;    
		mem[   497] = 11'd27;    
		mem[   498] = 11'd23;    
		mem[   499] = 11'd52;    
		mem[   500] = 11'd47;    
		mem[   501] = 11'd51;    
		mem[   502] = 11'd44;    
		mem[   503] = 11'd28;    
		mem[   504] = 11'd22;    
		mem[   505] = 11'd53;    
		mem[   506] = 11'd47;    
		mem[   507] = 11'd50;    
		mem[   508] = 11'd46;    
		mem[   509] = 11'd26;    
		mem[   510] = 11'd23;    
		mem[   511] = 11'd52;    
		mem[   512] = 11'd47;    
		mem[   513] = 11'd51;    
		mem[   514] = 11'd49;    
		mem[   515] = 11'd26;    
		mem[   516] = 11'd22;    
		mem[   517] = 11'd25;    
		mem[   518] = 11'd24;    
		mem[   519] = 11'd25;    
		mem[   520] = 11'd23;    
		mem[   521] = 11'd25;    
		mem[   522] = 11'd24;    
		mem[   523] = 11'd25;    
		mem[   524] = 11'd24;    
		mem[   525] = 11'd24;    
		mem[   526] = 11'd25;    
		mem[   527] = 11'd24;    
		mem[   528] = 11'd25;    
		mem[   529] = 11'd24;    
		mem[   530] = 11'd25;    
		mem[   531] = 11'd24;    
		mem[   532] = 11'd25;    
		mem[   533] = 11'd24;    
		mem[   534] = 11'd25;    
		mem[   535] = 11'd24;    
		mem[   536] = 11'd25;    
		mem[   537] = 11'd24;    
		mem[   538] = 11'd25;    
		mem[   539] = 11'd24;    
		mem[   540] = 11'd25;    
		mem[   541] = 11'd24;    
		mem[   542] = 11'd25;    
		mem[   543] = 11'd23;    
		mem[   544] = 11'd26;    
		mem[   545] = 11'd98;    
		mem[   546] = 11'd50;    
		mem[   547] = 11'd25;    
		mem[   548] = 11'd24;    
		mem[   549] = 11'd47;    
		mem[   550] = 11'd50;    
		mem[   551] = 11'd50;    
		mem[   552] = 11'd25;    
		mem[   553] = 11'd24;    
		mem[   554] = 11'd47;    
		mem[   555] = 11'd50;    
		mem[   556] = 11'd50;    
		mem[   557] = 11'd24;    
		mem[   558] = 11'd25;    
		mem[   559] = 11'd46;    
		mem[   560] = 11'd50;    
		mem[   561] = 11'd50;    
		mem[   562] = 11'd25;    
		mem[   563] = 11'd24;    
		mem[   564] = 11'd47;    
		mem[   565] = 11'd50;    
		mem[   566] = 11'd50;    
		mem[   567] = 11'd25;    
		mem[   568] = 11'd24;    
		mem[   569] = 11'd47;    
		mem[   570] = 11'd50;    
		mem[   571] = 11'd49;    
		mem[   572] = 11'd25;    
		mem[   573] = 11'd24;    
		mem[   574] = 11'd48;    
		mem[   575] = 11'd50;    
		mem[   576] = 11'd49;    
		mem[   577] = 11'd25;    
		mem[   578] = 11'd24;    
		mem[   579] = 11'd47;    
		mem[   580] = 11'd49;    
		mem[   581] = 11'd24;    
		mem[   582] = 11'd25;    
		mem[   583] = 11'd25;    
		mem[   584] = 11'd24;    
		mem[   585] = 11'd25;    
		mem[   586] = 11'd24;    
		mem[   587] = 11'd26;    
		mem[   588] = 11'd23;    
		mem[   589] = 11'd25;    
		mem[   590] = 11'd24;    
		mem[   591] = 11'd25;    
		mem[   592] = 11'd24;    
		mem[   593] = 11'd75;    
		mem[   594] = 11'd22;    
		mem[   595] = 11'd49;    
		mem[   596] = 11'd24;    
		mem[   597] = 11'd76;    
		mem[   598] = 11'd48;    
		mem[   599] = 11'd27;    
		mem[   600] = 11'd9;    
		mem[   601] = 11'd15;    
		mem[   602] = 11'd46;    
		mem[   603] = 11'd50;    
		mem[   604] = 11'd51;    
		mem[   605] = 11'd22;    
		mem[   606] = 11'd24;    
		mem[   607] = 11'd51;    
		mem[   608] = 11'd46;    
		mem[   609] = 11'd52;    
		mem[   610] = 11'd37;    
		mem[   611] = 11'd8;    
		mem[   612] = 11'd53;    
		mem[   613] = 11'd24;    
		mem[   614] = 11'd72;    
		mem[   615] = 11'd25;    
		mem[   616] = 11'd75;    
		mem[   617] = 11'd20;    
		mem[   618] = 11'd26;    
		mem[   619] = 11'd46;    
		mem[   620] = 11'd14;    
		mem[   621] = 11'd38;    
		mem[   622] = 11'd50;    
		mem[   623] = 11'd50;    
		mem[   624] = 11'd24;    
		mem[   625] = 11'd24;    
		mem[   626] = 11'd49;    
		mem[   627] = 11'd48;    
		mem[   628] = 11'd51;    
		mem[   629] = 11'd47;    
		mem[   630] = 11'd48;    
		mem[   631] = 11'd50;    
		mem[   632] = 11'd24;    
		mem[   633] = 11'd25;    
		mem[   634] = 11'd25;    
		mem[   635] = 11'd24;    
		mem[   636] = 11'd25;    
		mem[   637] = 11'd24;    
		mem[   638] = 11'd25;    
		mem[   639] = 11'd24;    
		mem[   640] = 11'd25;    
		mem[   641] = 11'd24;    
		mem[   642] = 11'd25;    
		mem[   643] = 11'd25;    
		mem[   644] = 11'd49;    
		mem[   645] = 11'd71;    
		mem[   646] = 11'd25;    
		mem[   647] = 11'd52;    
		mem[   648] = 11'd24;    
		mem[   649] = 11'd71;    
		mem[   650] = 11'd24;    
		mem[   651] = 11'd75;    
		mem[   652] = 11'd50;    
		mem[   653] = 11'd23;    
		mem[   654] = 11'd24;    
		mem[   655] = 11'd50;    
		mem[   656] = 11'd46;    
		mem[   657] = 11'd52;    
		mem[   658] = 11'd24;    
		mem[   659] = 11'd87;    
		mem[   660] = 11'd65;    
		mem[   661] = 11'd23;    
		mem[   662] = 11'd86;    
		mem[   663] = 11'd65;    
		mem[   664] = 11'd23;    
		mem[   665] = 11'd86;    
		mem[   666] = 11'd66;    
		mem[   667] = 11'd22;    
		mem[   668] = 11'd86;    
		mem[   669] = 11'd66;    
		mem[   670] = 11'd22;    
		mem[   671] = 11'd247;    
		mem[   672] = 11'd264;    
		mem[   673] = 11'd21;    
		mem[   674] = 11'd82;    
		mem[   675] = 11'd62;    
		mem[   676] = 11'd21;    
		mem[   677] = 11'd82;    
		mem[   678] = 11'd63;    
		mem[   679] = 11'd21;    
		mem[   680] = 11'd80;    
		mem[   681] = 11'd63;    
		mem[   682] = 11'd21;    
		mem[   683] = 11'd79;    
		mem[   684] = 11'd63;    
		mem[   685] = 11'd21;    
		mem[   686] = 11'd80;    
		mem[   687] = 11'd62;    
		mem[   688] = 11'd21;    
		mem[   689] = 11'd81;    
		mem[   690] = 11'd61;    
		mem[   691] = 11'd22;    
		mem[   692] = 11'd81;    
		mem[   693] = 11'd61;    
		mem[   694] = 11'd21;    
		mem[   695] = 11'd82;    
		mem[   696] = 11'd61;    
		mem[   697] = 11'd21;    
		mem[   698] = 11'd251;    
		mem[   699] = 11'd202;    
		mem[   700] = 11'd67;    
		mem[   701] = 11'd30;    
		mem[   702] = 11'd33;    
		mem[   703] = 11'd68;    
		mem[   704] = 11'd61;    
		mem[   705] = 11'd69;    
		mem[   706] = 11'd61;    
		mem[   707] = 11'd70;    
		mem[   708] = 11'd32;    
		mem[   709] = 11'd15;    
		mem[   710] = 11'd80;    
		mem[   711] = 11'd33;    
		mem[   712] = 11'd98;    
		mem[   713] = 11'd28;    
		mem[   714] = 11'd29;    
		mem[   715] = 11'd63;    
		mem[   716] = 11'd31;    
		mem[   717] = 11'd94;    
		mem[   718] = 11'd28;    
		mem[   719] = 11'd29;    
		mem[   720] = 11'd63;    
		mem[   721] = 11'd31;    
		mem[   722] = 11'd28;    
		mem[   723] = 11'd66;    
		mem[   724] = 11'd28;    
		mem[   725] = 11'd29;    
		mem[   726] = 11'd63;    
		mem[   727] = 11'd31;    
		mem[   728] = 11'd94;    
		mem[   729] = 11'd28;    
		mem[   730] = 11'd30;    
		mem[   731] = 11'd62;    
		mem[   732] = 11'd31;    
		mem[   733] = 11'd28;    
		mem[   734] = 11'd37;    
		mem[   735] = 11'd29;    
		mem[   736] = 11'd28;    
		mem[   737] = 11'd29;    
		mem[   738] = 11'd63;    
		mem[   739] = 11'd31;    
		mem[   740] = 11'd29;    
		mem[   741] = 11'd36;    
		mem[   742] = 11'd29;    
		mem[   743] = 11'd28;    
		mem[   744] = 11'd30;    
		mem[   745] = 11'd62;    
		mem[   746] = 11'd31;    
		mem[   747] = 11'd29;    
		mem[   748] = 11'd35;    
		mem[   749] = 11'd30;    
		mem[   750] = 11'd29;    
		mem[   751] = 11'd29;    
		mem[   752] = 11'd62;    
		mem[   753] = 11'd31;    
		mem[   754] = 11'd29;    
		mem[   755] = 11'd35;    
		mem[   756] = 11'd30;    
		mem[   757] = 11'd29;    
		mem[   758] = 11'd29;    
		mem[   759] = 11'd35;    
		mem[   760] = 11'd28;    
		mem[   761] = 11'd30;    
		mem[   762] = 11'd30;    
		mem[   763] = 11'd34;    
		mem[   764] = 11'd29;    
		mem[   765] = 11'd30;    
		mem[   766] = 11'd17;    
		mem[   767] = 11'd13;    
		mem[   768] = 11'd62;    
		mem[   769] = 11'd31;    
		mem[   770] = 11'd17;    
		mem[   771] = 11'd12;    
		mem[   772] = 11'd31;    
		mem[   773] = 11'd31;    
		mem[   774] = 11'd31;    
		mem[   775] = 11'd31;    
		mem[   776] = 11'd31;    
		mem[   777] = 11'd30;    
		mem[   778] = 11'd31;    
		mem[   779] = 11'd30;    
		mem[   780] = 11'd32;    
		mem[   781] = 11'd30;    
		mem[   782] = 11'd31;    
		mem[   783] = 11'd30;    
		mem[   784] = 11'd31;    
		mem[   785] = 11'd30;    
		mem[   786] = 11'd31;    
		mem[   787] = 11'd30;    
		mem[   788] = 11'd32;    
		mem[   789] = 11'd29;    
		mem[   790] = 11'd32;    
		mem[   791] = 11'd30;    
		mem[   792] = 11'd31;    
		mem[   793] = 11'd30;    
		mem[   794] = 11'd31;    
		mem[   795] = 11'd30;    
		mem[   796] = 11'd32;    
		mem[   797] = 11'd32;    
		mem[   798] = 11'd33;    
		mem[   799] = 11'd32;    
		mem[   800] = 11'd33;    
		mem[   801] = 11'd32;    
		mem[   802] = 11'd33;    
		mem[   803] = 11'd32;    
		mem[   804] = 11'd33;    
		mem[   805] = 11'd32;    
		mem[   806] = 11'd33;    
		mem[   807] = 11'd32;    
		mem[   808] = 11'd33;    
		mem[   809] = 11'd32;    
		mem[   810] = 11'd33;    
		mem[   811] = 11'd32;    
		mem[   812] = 11'd33;    
		mem[   813] = 11'd32;    
		mem[   814] = 11'd33;    
		mem[   815] = 11'd32;    
		mem[   816] = 11'd33;    
		mem[   817] = 11'd32;    
		mem[   818] = 11'd33;    
		mem[   819] = 11'd30;    
		mem[   820] = 11'd31;    
		mem[   821] = 11'd30;    
		mem[   822] = 11'd31;    
		mem[   823] = 11'd30;    
		mem[   824] = 11'd32;    
		mem[   825] = 11'd30;    
		mem[   826] = 11'd31;    
		mem[   827] = 11'd30;    
		mem[   828] = 11'd31;    
		mem[   829] = 11'd30;    
		mem[   830] = 11'd31;    
		mem[   831] = 11'd30;    
		mem[   832] = 11'd32;    
		mem[   833] = 11'd30;    
		mem[   834] = 11'd31;    
		mem[   835] = 11'd30;    
		mem[   836] = 11'd31;    
		mem[   837] = 11'd30;    
		mem[   838] = 11'd32;    
		mem[   839] = 11'd30;    
		mem[   840] = 11'd31;    
		mem[   841] = 11'd30;    
		mem[   842] = 11'd64;    
		mem[   843] = 11'd27;    
		mem[   844] = 11'd92;    
		mem[   845] = 11'd31;    
		mem[   846] = 11'd94;    
		mem[   847] = 11'd28;    
		mem[   848] = 11'd92;    
		mem[   849] = 11'd31;    
		mem[   850] = 11'd94;    
		mem[   851] = 11'd28;    
		mem[   852] = 11'd92;    
		mem[   853] = 11'd31;    
		mem[   854] = 11'd94;    
		mem[   855] = 11'd28;    
		mem[   856] = 11'd30;    
		mem[   857] = 11'd63;    
		mem[   858] = 11'd30;    
		mem[   859] = 11'd94;    
		mem[   860] = 11'd29;    
		mem[   861] = 11'd28;    
		mem[   862] = 11'd64;    
		mem[   863] = 11'd30;    
		mem[   864] = 11'd29;    
		mem[   865] = 11'd65;    
		mem[   866] = 11'd29;    
		mem[   867] = 11'd29;    
		mem[   868] = 11'd63;    
		mem[   869] = 11'd31;    
		mem[   870] = 11'd28;    
		mem[   871] = 11'd63;    
		mem[   872] = 11'd31;    
		mem[   873] = 11'd31;    
		mem[   874] = 11'd31;    
		mem[   875] = 11'd30;    
		mem[   876] = 11'd32;    
		mem[   877] = 11'd30;    
		mem[   878] = 11'd31;    
		mem[   879] = 11'd30;    
		mem[   880] = 11'd31;    
		mem[   881] = 11'd30;    
		mem[   882] = 11'd32;    
		mem[   883] = 11'd29;    
		mem[   884] = 11'd32;    
		mem[   885] = 11'd30;    
		mem[   886] = 11'd31;    
		mem[   887] = 11'd30;    
		mem[   888] = 11'd31;    
		mem[   889] = 11'd30;    
		mem[   890] = 11'd31;    
		mem[   891] = 11'd30;    
		mem[   892] = 11'd32;    
		mem[   893] = 11'd30;    
		mem[   894] = 11'd67;    
		mem[   895] = 11'd63;    
		mem[   896] = 11'd36;    
		mem[   897] = 11'd12;    
		mem[   898] = 11'd19;    
		mem[   899] = 11'd62;    
		mem[   900] = 11'd65;    
		mem[   901] = 11'd67;    
		mem[   902] = 11'd30;    
		mem[   903] = 11'd32;    
		mem[   904] = 11'd67;    
		mem[   905] = 11'd36;    
		mem[   906] = 11'd26;    
		mem[   907] = 11'd69;    
		mem[   908] = 11'd49;    
		mem[   909] = 11'd78;    
		mem[   910] = 11'd30;    
		mem[   911] = 11'd15;    
		mem[   912] = 11'd77;    
		mem[   913] = 11'd36;    
		mem[   914] = 11'd10;    
		mem[   915] = 11'd12;    
		mem[   916] = 11'd66;    
		mem[   917] = 11'd30;    
		mem[   918] = 11'd14;    
		mem[   919] = 11'd77;    
		mem[   920] = 11'd36;    
		mem[   921] = 11'd11;    
		mem[   922] = 11'd11;    
		mem[   923] = 11'd66;    
		mem[   924] = 11'd30;    
		mem[   925] = 11'd14;    
		mem[   926] = 11'd77;    
		mem[   927] = 11'd36;    
		mem[   928] = 11'd11;    
		mem[   929] = 11'd11;    
		mem[   930] = 11'd65;    
		mem[   931] = 11'd31;    
		mem[   932] = 11'd15;    
		mem[   933] = 11'd12;    
		mem[   934] = 11'd64;    
		mem[   935] = 11'd36;    
		mem[   936] = 11'd23;    
		mem[   937] = 11'd65;    
		mem[   938] = 11'd30;    
		mem[   939] = 11'd15;    
		mem[   940] = 11'd12;    
		mem[   941] = 11'd36;    
		mem[   942] = 11'd28;    
		mem[   943] = 11'd36;    
		mem[   944] = 11'd23;    
		mem[   945] = 11'd64;    
		mem[   946] = 11'd14;    
		mem[   947] = 11'd17;    
		mem[   948] = 11'd15;    
		mem[   949] = 11'd12;    
		mem[   950] = 11'd36;    
		mem[   951] = 11'd28;    
		mem[   952] = 11'd36;    
		mem[   953] = 11'd23;    
		mem[   954] = 11'd64;    
		mem[   955] = 11'd31;    
		mem[   956] = 11'd16;    
		mem[   957] = 11'd11;    
		mem[   958] = 11'd36;    
		mem[   959] = 11'd28;    
		mem[   960] = 11'd36;    
		mem[   961] = 11'd23;    
		mem[   962] = 11'd65;    
		mem[   963] = 11'd30;    
		mem[   964] = 11'd27;    
		mem[   965] = 11'd35;    
		mem[   966] = 11'd29;    
		mem[   967] = 11'd33;    
		mem[   968] = 11'd27;    
		mem[   969] = 11'd31;    
		mem[   970] = 11'd32;    
		mem[   971] = 11'd31;    
		mem[   972] = 11'd28;    
		mem[   973] = 11'd34;    
		mem[   974] = 11'd29;    
		mem[   975] = 11'd33;    
		mem[   976] = 11'd26;    
		mem[   977] = 11'd62;    
		mem[   978] = 11'd31;    
		mem[   979] = 11'd31;    
		mem[   980] = 11'd31;    
		mem[   981] = 11'd30;    
		mem[   982] = 11'd32;    
		mem[   983] = 11'd30;    
		mem[   984] = 11'd31;    
		mem[   985] = 11'd30;    
		mem[   986] = 11'd32;    
		mem[   987] = 11'd30;    
		mem[   988] = 11'd31;    
		mem[   989] = 11'd30;    
		mem[   990] = 11'd31;    
		mem[   991] = 11'd30;    
		mem[   992] = 11'd31;    
		mem[   993] = 11'd30;    
		mem[   994] = 11'd31;    
		mem[   995] = 11'd30;    
		mem[   996] = 11'd32;    
		mem[   997] = 11'd30;    
		mem[   998] = 11'd31;    
		mem[   999] = 11'd33;    
		mem[  1000] = 11'd39;    
		mem[  1001] = 11'd38;    
		mem[  1002] = 11'd40;    
		mem[  1003] = 11'd38;    
		mem[  1004] = 11'd40;    
		mem[  1005] = 11'd38;    
		mem[  1006] = 11'd39;    
		mem[  1007] = 11'd38;    
		mem[  1008] = 11'd40;    
		mem[  1009] = 11'd38;    
		mem[  1010] = 11'd39;    
		mem[  1011] = 11'd39;    
		mem[  1012] = 11'd39;    
		mem[  1013] = 11'd38;    
		mem[  1014] = 11'd40;    
		mem[  1015] = 11'd38;    
		mem[  1016] = 11'd40;    
		mem[  1017] = 11'd38;    
		mem[  1018] = 11'd38;    
		mem[  1019] = 11'd36;    
		mem[  1020] = 11'd37;    
		mem[  1021] = 11'd36;    
		mem[  1022] = 11'd37;    
		mem[  1023] = 11'd36;    
		mem[  1024] = 11'd37;    
		mem[  1025] = 11'd36;    
		mem[  1026] = 11'd38;    
		mem[  1027] = 11'd35;    
		mem[  1028] = 11'd38;    
		mem[  1029] = 11'd36;    
		mem[  1030] = 11'd37;    
		mem[  1031] = 11'd36;    
		mem[  1032] = 11'd37;    
		mem[  1033] = 11'd36;    
		mem[  1034] = 11'd37;    
		mem[  1035] = 11'd36;    
		mem[  1036] = 11'd38;    
		mem[  1037] = 11'd35;    
		mem[  1038] = 11'd37;    
		mem[  1039] = 11'd76;    
		mem[  1040] = 11'd102;    
		mem[  1041] = 11'd22;    
		mem[  1042] = 11'd55;    
		mem[  1043] = 11'd74;    
		mem[  1044] = 11'd75;    
		mem[  1045] = 11'd41;    
		mem[  1046] = 11'd106;    
		mem[  1047] = 11'd72;    
		mem[  1048] = 11'd37;    
		mem[  1049] = 11'd35;    
		mem[  1050] = 11'd83;    
		mem[  1051] = 11'd19;    
		mem[  1052] = 11'd19;    
		mem[  1053] = 11'd40;    
		mem[  1054] = 11'd46;    
		mem[  1055] = 11'd37;    
		mem[  1056] = 11'd85;    
		mem[  1057] = 11'd20;    
		mem[  1058] = 11'd18;    
		mem[  1059] = 11'd40;    
		mem[  1060] = 11'd46;    
		mem[  1061] = 11'd37;    
		mem[  1062] = 11'd85;    
		mem[  1063] = 11'd18;    
		mem[  1064] = 11'd20;    
		mem[  1065] = 11'd40;    
		mem[  1066] = 11'd45;    
		mem[  1067] = 11'd38;    
		mem[  1068] = 11'd41;    
		mem[  1069] = 11'd41;    
		mem[  1070] = 11'd41;    
		mem[  1071] = 11'd41;    
		mem[  1072] = 11'd41;    
		mem[  1073] = 11'd41;    
		mem[  1074] = 11'd41;    
		mem[  1075] = 11'd41;    
		mem[  1076] = 11'd41;    
		mem[  1077] = 11'd40;    
		mem[  1078] = 11'd42;    
		mem[  1079] = 11'd40;    
		mem[  1080] = 11'd42;    
		mem[  1081] = 11'd40;    
		mem[  1082] = 11'd42;    
		mem[  1083] = 11'd40;    
		mem[  1084] = 11'd42;    
		mem[  1085] = 11'd38;    
		mem[  1086] = 11'd64;    
		mem[  1087] = 11'd57;    
		mem[  1088] = 11'd66;    
		mem[  1089] = 11'd57;    
		mem[  1090] = 11'd65;    
		mem[  1091] = 11'd57;    
		mem[  1092] = 11'd66;    
		mem[  1093] = 11'd57;    
		mem[  1094] = 11'd65;    
		mem[  1095] = 11'd58;    
		mem[  1096] = 11'd65;    
		mem[  1097] = 11'd58;    
		mem[  1098] = 11'd64;    
		mem[  1099] = 11'd58;    
		mem[  1100] = 11'd65;    
		mem[  1101] = 11'd58;    
		mem[  1102] = 11'd64;    
		mem[  1103] = 11'd58;    
		mem[  1104] = 11'd65;    
		mem[  1105] = 11'd58;    
		mem[  1106] = 11'd64;    
		mem[  1107] = 11'd58;    
		mem[  1108] = 11'd65;    
		mem[  1109] = 11'd24;    
		mem[  1110] = 11'd33;    
		mem[  1111] = 11'd114;    
		mem[  1112] = 11'd91;    
		mem[  1113] = 11'd31;    
		mem[  1114] = 11'd121;    
		mem[  1115] = 11'd93;    
		mem[  1116] = 11'd31;    
		mem[  1117] = 11'd122;    
		mem[  1118] = 11'd92;    
		mem[  1119] = 11'd35;    
		mem[  1120] = 11'd62;    
		mem[  1121] = 11'd34;    
		mem[  1122] = 11'd27;    
		mem[  1123] = 11'd63;    
		mem[  1124] = 11'd29;    
		mem[  1125] = 11'd31;    
		mem[  1126] = 11'd62;    
		mem[  1127] = 11'd60;    
		mem[  1128] = 11'd63;    
		mem[  1129] = 11'd30;    
		mem[  1130] = 11'd30;    
		mem[  1131] = 11'd62;    
		mem[  1132] = 11'd34;    
		mem[  1133] = 11'd26;    
		mem[  1134] = 11'd63;    
		mem[  1135] = 11'd30;    
		mem[  1136] = 11'd28;    
		mem[  1137] = 11'd62;    
		mem[  1138] = 11'd31;    
		mem[  1139] = 11'd31;    
		mem[  1140] = 11'd32;    
		mem[  1141] = 11'd30;    
		mem[  1142] = 11'd31;    
		mem[  1143] = 11'd30;    
		mem[  1144] = 11'd32;    
		mem[  1145] = 11'd30;    
		mem[  1146] = 11'd31;    
		mem[  1147] = 11'd30;    
		mem[  1148] = 11'd32;    
		mem[  1149] = 11'd29;    
		mem[  1150] = 11'd32;    
		mem[  1151] = 11'd29;    
		mem[  1152] = 11'd32;    
		mem[  1153] = 11'd30;    
		mem[  1154] = 11'd31;    
		mem[  1155] = 11'd30;    
		mem[  1156] = 11'd31;    
		mem[  1157] = 11'd30;    
		mem[  1158] = 11'd32;    
		mem[  1159] = 11'd29;    
		mem[  1160] = 11'd32;    
		mem[  1161] = 11'd30;    
		mem[  1162] = 11'd31;    
		mem[  1163] = 11'd30;    
		mem[  1164] = 11'd31;    
		mem[  1165] = 11'd30;    
		mem[  1166] = 11'd31;    
		mem[  1167] = 11'd30;    
		mem[  1168] = 11'd32;    
		mem[  1169] = 11'd30;    
		mem[  1170] = 11'd31;    
		mem[  1171] = 11'd30;    
		mem[  1172] = 11'd31;    
		mem[  1173] = 11'd30;    
		mem[  1174] = 11'd31;    
		mem[  1175] = 11'd30;    
		mem[  1176] = 11'd32;    
		mem[  1177] = 11'd30;    
		mem[  1178] = 11'd31;    
		mem[  1179] = 11'd30;    
		mem[  1180] = 11'd31;    
		mem[  1181] = 11'd30;    
		mem[  1182] = 11'd31;    
		mem[  1183] = 11'd30;    
		mem[  1184] = 11'd31;    
		mem[  1185] = 11'd31;    
		mem[  1186] = 11'd30;    
		mem[  1187] = 11'd31;    
		mem[  1188] = 11'd31;    
		mem[  1189] = 11'd30;    
		mem[  1190] = 11'd31;    
		mem[  1191] = 11'd30;    
		mem[  1192] = 11'd31;    
		mem[  1193] = 11'd31;    
		mem[  1194] = 11'd31;    
		mem[  1195] = 11'd30;    
		mem[  1196] = 11'd31;    
		mem[  1197] = 11'd30;    
		mem[  1198] = 11'd31;    
		mem[  1199] = 11'd31;    
		mem[  1200] = 11'd31;    
		mem[  1201] = 11'd30;    
		mem[  1202] = 11'd31;    
		mem[  1203] = 11'd30;    
		mem[  1204] = 11'd31;    
		mem[  1205] = 11'd30;    
		mem[  1206] = 11'd72;    
		mem[  1207] = 11'd81;    
		mem[  1208] = 11'd79;    
		mem[  1209] = 11'd57;    
		mem[  1210] = 11'd58;    
		mem[  1211] = 11'd39;    
		mem[  1212] = 11'd78;    
		mem[  1213] = 11'd35;    
		mem[  1214] = 11'd38;    
		mem[  1215] = 11'd83;    
		mem[  1216] = 11'd35;    
		mem[  1217] = 11'd39;    
		mem[  1218] = 11'd43;    
		mem[  1219] = 11'd35;    
		mem[  1220] = 11'd74;    
		mem[  1221] = 11'd39;    
		mem[  1222] = 11'd17;    
		mem[  1223] = 11'd88;    
		mem[  1224] = 11'd35;    
		mem[  1225] = 11'd37;    
		mem[  1226] = 11'd75;    
		mem[  1227] = 11'd76;    
		mem[  1228] = 11'd68;    
		mem[  1229] = 11'd38;    
		mem[  1230] = 11'd40;    
		mem[  1231] = 11'd32;    
		mem[  1232] = 11'd38;    
		mem[  1233] = 11'd41;    
		mem[  1234] = 11'd34;    
		mem[  1235] = 11'd38;    
		mem[  1236] = 11'd34;    
		mem[  1237] = 11'd37;    
		mem[  1238] = 11'd36;    
		mem[  1239] = 11'd37;    
		mem[  1240] = 11'd36;    
		mem[  1241] = 11'd37;    
		mem[  1242] = 11'd36;    
		mem[  1243] = 11'd37;    
		mem[  1244] = 11'd36;    
		mem[  1245] = 11'd37;    
		mem[  1246] = 11'd37;    
		mem[  1247] = 11'd36;    
		mem[  1248] = 11'd37;    
		mem[  1249] = 11'd37;    
		mem[  1250] = 11'd36;    
		mem[  1251] = 11'd37;    
		mem[  1252] = 11'd36;    
		mem[  1253] = 11'd37;    
		mem[  1254] = 11'd35;    
		mem[  1255] = 11'd77;    
		mem[  1256] = 11'd74;    
		mem[  1257] = 11'd40;    
		mem[  1258] = 11'd103;    
		mem[  1259] = 11'd73;    
		mem[  1260] = 11'd19;    
		mem[  1261] = 11'd55;    
		mem[  1262] = 11'd39;    
		mem[  1263] = 11'd16;    
		mem[  1264] = 11'd61;    
		mem[  1265] = 11'd7;    
		mem[  1266] = 11'd23;    
		mem[  1267] = 11'd76;    
		mem[  1268] = 11'd73;    
		mem[  1269] = 11'd14;    
		mem[  1270] = 11'd20;    
		mem[  1271] = 11'd20;    
		mem[  1272] = 11'd13;    
		mem[  1273] = 11'd76;    
		mem[  1274] = 11'd73;    
		mem[  1275] = 11'd74;    
		mem[  1276] = 11'd40;    
		mem[  1277] = 11'd16;    
		mem[  1278] = 11'd58;    
		mem[  1279] = 11'd12;    
		mem[  1280] = 11'd20;    
		mem[  1281] = 11'd76;    
		mem[  1282] = 11'd73;    
		mem[  1283] = 11'd14;    
		mem[  1284] = 11'd41;    
		mem[  1285] = 11'd13;    
		mem[  1286] = 11'd77;    
		mem[  1287] = 11'd38;    
		mem[  1288] = 11'd34;    
		mem[  1289] = 11'd38;    
		mem[  1290] = 11'd35;    
		mem[  1291] = 11'd37;    
		mem[  1292] = 11'd36;    
		mem[  1293] = 11'd37;    
		mem[  1294] = 11'd36;    
		mem[  1295] = 11'd39;    
		mem[  1296] = 11'd33;    
		mem[  1297] = 11'd42;    
		mem[  1298] = 11'd30;    
		mem[  1299] = 11'd78;    
		mem[  1300] = 11'd34;    
		mem[  1301] = 11'd38;    
		mem[  1302] = 11'd34;    
		mem[  1303] = 11'd24;    
		mem[  1304] = 11'd88;    
		mem[  1305] = 11'd72;    
		mem[  1306] = 11'd19;    
		mem[  1307] = 11'd56;    
		mem[  1308] = 11'd37;    
		mem[  1309] = 11'd35;    
		mem[  1310] = 11'd37;    
		mem[  1311] = 11'd34;    
		mem[  1312] = 11'd76;    
		mem[  1313] = 11'd73;    
		mem[  1314] = 11'd74;    
		mem[  1315] = 11'd38;    
		mem[  1316] = 11'd32;    
		mem[  1317] = 11'd40;    
		mem[  1318] = 11'd33;    
		mem[  1319] = 11'd40;    
		mem[  1320] = 11'd36;    
		mem[  1321] = 11'd73;    
		mem[  1322] = 11'd33;    
		mem[  1323] = 11'd39;    
		mem[  1324] = 11'd40;    
		mem[  1325] = 11'd17;    
		mem[  1326] = 11'd15;    
		mem[  1327] = 11'd42;    
		mem[  1328] = 11'd32;    
		mem[  1329] = 11'd59;    
		mem[  1330] = 11'd14;    
		mem[  1331] = 11'd37;    
		mem[  1332] = 11'd37;    
		mem[  1333] = 11'd37;    
		mem[  1334] = 11'd36;    
		mem[  1335] = 11'd38;    
		mem[  1336] = 11'd36;    
		mem[  1337] = 11'd37;    
		mem[  1338] = 11'd36;    
		mem[  1339] = 11'd75;    
		mem[  1340] = 11'd71;    
		mem[  1341] = 11'd20;    
		mem[  1342] = 11'd56;    
		mem[  1343] = 11'd34;    
		mem[  1344] = 11'd38;    
		mem[  1345] = 11'd30;    
		mem[  1346] = 11'd25;    
		mem[  1347] = 11'd87;    
		mem[  1348] = 11'd62;    
		mem[  1349] = 11'd16;    
		mem[  1350] = 11'd73;    
		mem[  1351] = 11'd73;    
		mem[  1352] = 11'd34;    
		mem[  1353] = 11'd36;    
		mem[  1354] = 11'd41;    
		mem[  1355] = 11'd70;    
		mem[  1356] = 11'd23;    
		mem[  1357] = 11'd87;    
		mem[  1358] = 11'd68;    
		mem[  1359] = 11'd22;    
		mem[  1360] = 11'd84;    
		mem[  1361] = 11'd68;    
		mem[  1362] = 11'd22;    
		mem[  1363] = 11'd85;    
		mem[  1364] = 11'd67;    
		mem[  1365] = 11'd23;    
		mem[  1366] = 11'd84;    
		mem[  1367] = 11'd430;    
		mem[  1368] = 11'd21;    
		mem[  1369] = 11'd80;    
		mem[  1370] = 11'd61;    
		mem[  1371] = 11'd20;    
		mem[  1372] = 11'd80;    
		mem[  1373] = 11'd61;    
		mem[  1374] = 11'd22;    
		mem[  1375] = 11'd81;    
		mem[  1376] = 11'd61;    
		mem[  1377] = 11'd21;    
		mem[  1378] = 11'd82;    
		mem[  1379] = 11'd62;    
		mem[  1380] = 11'd21;    
		mem[  1381] = 11'd80;    
		mem[  1382] = 11'd62;    
		mem[  1383] = 11'd22;    
		mem[  1384] = 11'd80;    
		mem[  1385] = 11'd63;    
		mem[  1386] = 11'd21;    
		mem[  1387] = 11'd80;    
		mem[  1388] = 11'd63;    
		mem[  1389] = 11'd21;    
		mem[  1390] = 11'd80;    
		mem[  1391] = 11'd62;    
		mem[  1392] = 11'd22;    
		mem[  1393] = 11'd250;    
		mem[  1394] = 11'd197;    
		mem[  1395] = 11'd97;    
		mem[  1396] = 11'd33;    
		mem[  1397] = 11'd100;    
		mem[  1398] = 11'd63;    
		mem[  1399] = 11'd52;    
		mem[  1400] = 11'd13;    
		mem[  1401] = 11'd64;    
		mem[  1402] = 11'd66;    
		mem[  1403] = 11'd67;    
		mem[  1404] = 11'd30;    
		mem[  1405] = 11'd33;    
		mem[  1406] = 11'd66;    
		mem[  1407] = 11'd61;    
		mem[  1408] = 11'd65;    
		mem[  1409] = 11'd25;    
		mem[  1410] = 11'd33;    
		mem[  1411] = 11'd63;    
		mem[  1412] = 11'd59;    
		mem[  1413] = 11'd65;    
		mem[  1414] = 11'd26;    
		mem[  1415] = 11'd32;    
		mem[  1416] = 11'd63;    
		mem[  1417] = 11'd59;    
		mem[  1418] = 11'd65;    
		mem[  1419] = 11'd26;    
		mem[  1420] = 11'd32;    
		mem[  1421] = 11'd63;    
		mem[  1422] = 11'd59;    
		mem[  1423] = 11'd64;    
		mem[  1424] = 11'd27;    
		mem[  1425] = 11'd32;    
		mem[  1426] = 11'd63;    
		mem[  1427] = 11'd59;    
		mem[  1428] = 11'd65;    
		mem[  1429] = 11'd26;    
		mem[  1430] = 11'd32;    
		mem[  1431] = 11'd63;    
		mem[  1432] = 11'd59;    
		mem[  1433] = 11'd64;    
		mem[  1434] = 11'd27;    
		mem[  1435] = 11'd32;    
		mem[  1436] = 11'd63;    
		mem[  1437] = 11'd34;    
		mem[  1438] = 11'd26;    
		mem[  1439] = 11'd63;    
		mem[  1440] = 11'd27;    
		mem[  1441] = 11'd32;    
		mem[  1442] = 11'd63;    
		mem[  1443] = 11'd34;    
		mem[  1444] = 11'd26;    
		mem[  1445] = 11'd64;    
		mem[  1446] = 11'd27;    
		mem[  1447] = 11'd31;    
		mem[  1448] = 11'd63;    
		mem[  1449] = 11'd33;    
		mem[  1450] = 11'd27;    
		mem[  1451] = 11'd63;    
		mem[  1452] = 11'd28;    
		mem[  1453] = 11'd32;    
		mem[  1454] = 11'd62;    
		mem[  1455] = 11'd62;    
		mem[  1456] = 11'd32;    
		mem[  1457] = 11'd28;    
		mem[  1458] = 11'd32;    
		mem[  1459] = 11'd29;    
		mem[  1460] = 11'd31;    
		mem[  1461] = 11'd30;    
		mem[  1462] = 11'd31;    
		mem[  1463] = 11'd30;    
		mem[  1464] = 11'd31;    
		mem[  1465] = 11'd31;    
		mem[  1466] = 11'd30;    
		mem[  1467] = 11'd31;    
		mem[  1468] = 11'd30;    
		mem[  1469] = 11'd31;    
		mem[  1470] = 11'd31;    
		mem[  1471] = 11'd31;    
		mem[  1472] = 11'd30;    
		mem[  1473] = 11'd31;    
		mem[  1474] = 11'd31;    
		mem[  1475] = 11'd30;    
		mem[  1476] = 11'd31;    
		mem[  1477] = 11'd31;    
		mem[  1478] = 11'd32;    
		mem[  1479] = 11'd32;    
		mem[  1480] = 11'd33;    
		mem[  1481] = 11'd32;    
		mem[  1482] = 11'd33;    
		mem[  1483] = 11'd32;    
		mem[  1484] = 11'd33;    
		mem[  1485] = 11'd32;    
		mem[  1486] = 11'd33;    
		mem[  1487] = 11'd32;    
		mem[  1488] = 11'd33;    
		mem[  1489] = 11'd32;    
		mem[  1490] = 11'd33;    
		mem[  1491] = 11'd32;    
		mem[  1492] = 11'd33;    
		mem[  1493] = 11'd32;    
		mem[  1494] = 11'd33;    
		mem[  1495] = 11'd32;    
		mem[  1496] = 11'd33;    
		mem[  1497] = 11'd32;    
		mem[  1498] = 11'd33;    
		mem[  1499] = 11'd32;    
		mem[  1500] = 11'd33;    
		mem[  1501] = 11'd30;    
		mem[  1502] = 11'd31;    
		mem[  1503] = 11'd30;    
		mem[  1504] = 11'd31;    
		mem[  1505] = 11'd30;    
		mem[  1506] = 11'd31;    
		mem[  1507] = 11'd30;    
		mem[  1508] = 11'd31;    
		mem[  1509] = 11'd30;    
		mem[  1510] = 11'd31;    
		mem[  1511] = 11'd31;    
		mem[  1512] = 11'd30;    
		mem[  1513] = 11'd31;    
		mem[  1514] = 11'd31;    
		mem[  1515] = 11'd30;    
		mem[  1516] = 11'd31;    
		mem[  1517] = 11'd30;    
		mem[  1518] = 11'd32;    
		mem[  1519] = 11'd30;    
		mem[  1520] = 11'd31;    
		mem[  1521] = 11'd30;    
		mem[  1522] = 11'd31;    
		mem[  1523] = 11'd30;    
		mem[  1524] = 11'd32;    
		mem[  1525] = 11'd27;    
		mem[  1526] = 11'd66;    
		mem[  1527] = 11'd25;    
		mem[  1528] = 11'd33;    
		mem[  1529] = 11'd64;    
		mem[  1530] = 11'd58;    
		mem[  1531] = 11'd66;    
		mem[  1532] = 11'd12;    
		mem[  1533] = 11'd13;    
		mem[  1534] = 11'd32;    
		mem[  1535] = 11'd64;    
		mem[  1536] = 11'd58;    
		mem[  1537] = 11'd66;    
		mem[  1538] = 11'd11;    
		mem[  1539] = 11'd14;    
		mem[  1540] = 11'd32;    
		mem[  1541] = 11'd64;    
		mem[  1542] = 11'd59;    
		mem[  1543] = 11'd65;    
		mem[  1544] = 11'd25;    
		mem[  1545] = 11'd32;    
		mem[  1546] = 11'd64;    
		mem[  1547] = 11'd58;    
		mem[  1548] = 11'd65;    
		mem[  1549] = 11'd26;    
		mem[  1550] = 11'd32;    
		mem[  1551] = 11'd64;    
		mem[  1552] = 11'd59;    
		mem[  1553] = 11'd64;    
		mem[  1554] = 11'd26;    
		mem[  1555] = 11'd32;    
		mem[  1556] = 11'd64;    
		mem[  1557] = 11'd61;    
		mem[  1558] = 11'd31;    
		mem[  1559] = 11'd30;    
		mem[  1560] = 11'd31;    
		mem[  1561] = 11'd30;    
		mem[  1562] = 11'd31;    
		mem[  1563] = 11'd30;    
		mem[  1564] = 11'd30;    
		mem[  1565] = 11'd31;    
		mem[  1566] = 11'd31;    
		mem[  1567] = 11'd30;    
		mem[  1568] = 11'd31;    
		mem[  1569] = 11'd30;    
		mem[  1570] = 11'd31;    
		mem[  1571] = 11'd31;    
		mem[  1572] = 11'd31;    
		mem[  1573] = 11'd30;    
		mem[  1574] = 11'd31;    
		mem[  1575] = 11'd30;    
		mem[  1576] = 11'd31;    
		mem[  1577] = 11'd31;    
		mem[  1578] = 11'd31;    
		mem[  1579] = 11'd31;    
		mem[  1580] = 11'd34;    
		mem[  1581] = 11'd96;    
		mem[  1582] = 11'd36;    
		mem[  1583] = 11'd62;    
		mem[  1584] = 11'd34;    
		mem[  1585] = 11'd29;    
		mem[  1586] = 11'd97;    
		mem[  1587] = 11'd24;    
		mem[  1588] = 11'd8;    
		mem[  1589] = 11'd32;    
		mem[  1590] = 11'd69;    
		mem[  1591] = 11'd63;    
		mem[  1592] = 11'd36;    
		mem[  1593] = 11'd13;    
		mem[  1594] = 11'd18;    
		mem[  1595] = 11'd62;    
		mem[  1596] = 11'd63;    
		mem[  1597] = 11'd62;    
		mem[  1598] = 11'd31;    
		mem[  1599] = 11'd31;    
		mem[  1600] = 11'd59;    
		mem[  1601] = 11'd62;    
		mem[  1602] = 11'd62;    
		mem[  1603] = 11'd31;    
		mem[  1604] = 11'd30;    
		mem[  1605] = 11'd60;    
		mem[  1606] = 11'd62;    
		mem[  1607] = 11'd62;    
		mem[  1608] = 11'd31;    
		mem[  1609] = 11'd31;    
		mem[  1610] = 11'd59;    
		mem[  1611] = 11'd62;    
		mem[  1612] = 11'd62;    
		mem[  1613] = 11'd31;    
		mem[  1614] = 11'd31;    
		mem[  1615] = 11'd59;    
		mem[  1616] = 11'd62;    
		mem[  1617] = 11'd62;    
		mem[  1618] = 11'd31;    
		mem[  1619] = 11'd31;    
		mem[  1620] = 11'd59;    
		mem[  1621] = 11'd62;    
		mem[  1622] = 11'd62;    
		mem[  1623] = 11'd31;    
		mem[  1624] = 11'd31;    
		mem[  1625] = 11'd59;    
		mem[  1626] = 11'd62;    
		mem[  1627] = 11'd62;    
		mem[  1628] = 11'd31;    
		mem[  1629] = 11'd31;    
		mem[  1630] = 11'd59;    
		mem[  1631] = 11'd62;    
		mem[  1632] = 11'd62;    
		mem[  1633] = 11'd31;    
		mem[  1634] = 11'd30;    
		mem[  1635] = 11'd60;    
		mem[  1636] = 11'd62;    
		mem[  1637] = 11'd62;    
		mem[  1638] = 11'd31;    
		mem[  1639] = 11'd31;    
		mem[  1640] = 11'd46;    
		mem[  1641] = 11'd12;    
		mem[  1642] = 11'd62;    
		mem[  1643] = 11'd31;    
		mem[  1644] = 11'd31;    
		mem[  1645] = 11'd31;    
		mem[  1646] = 11'd30;    
		mem[  1647] = 11'd32;    
		mem[  1648] = 11'd30;    
		mem[  1649] = 11'd31;    
		mem[  1650] = 11'd30;    
		mem[  1651] = 11'd31;    
		mem[  1652] = 11'd30;    
		mem[  1653] = 11'd32;    
		mem[  1654] = 11'd30;    
		mem[  1655] = 11'd31;    
		mem[  1656] = 11'd30;    
		mem[  1657] = 11'd31;    
		mem[  1658] = 11'd30;    
		mem[  1659] = 11'd32;    
		mem[  1660] = 11'd29;    
		mem[  1661] = 11'd31;    
		mem[  1662] = 11'd31;    
		mem[  1663] = 11'd31;    
		mem[  1664] = 11'd36;    
		mem[  1665] = 11'd39;    
		mem[  1666] = 11'd38;    
		mem[  1667] = 11'd40;    
		mem[  1668] = 11'd38;    
		mem[  1669] = 11'd40;    
		mem[  1670] = 11'd38;    
		mem[  1671] = 11'd39;    
		mem[  1672] = 11'd38;    
		mem[  1673] = 11'd40;    
		mem[  1674] = 11'd38;    
		mem[  1675] = 11'd40;    
		mem[  1676] = 11'd38;    
		mem[  1677] = 11'd39;    
		mem[  1678] = 11'd38;    
		mem[  1679] = 11'd40;    
		mem[  1680] = 11'd38;    
		mem[  1681] = 11'd39;    
		mem[  1682] = 11'd39;    
		mem[  1683] = 11'd37;    
		mem[  1684] = 11'd36;    
		mem[  1685] = 11'd37;    
		mem[  1686] = 11'd36;    
		mem[  1687] = 11'd37;    
		mem[  1688] = 11'd36;    
		mem[  1689] = 11'd38;    
		mem[  1690] = 11'd35;    
		mem[  1691] = 11'd38;    
		mem[  1692] = 11'd36;    
		mem[  1693] = 11'd37;    
		mem[  1694] = 11'd36;    
		mem[  1695] = 11'd37;    
		mem[  1696] = 11'd36;    
		mem[  1697] = 11'd37;    
		mem[  1698] = 11'd36;    
		mem[  1699] = 11'd37;    
		mem[  1700] = 11'd36;    
		mem[  1701] = 11'd37;    
		mem[  1702] = 11'd36;    
		mem[  1703] = 11'd75;    
		mem[  1704] = 11'd75;    
		mem[  1705] = 11'd14;    
		mem[  1706] = 11'd14;    
		mem[  1707] = 11'd39;    
		mem[  1708] = 11'd79;    
		mem[  1709] = 11'd32;    
		mem[  1710] = 11'd80;    
		mem[  1711] = 11'd15;    
		mem[  1712] = 11'd18;    
		mem[  1713] = 11'd72;    
		mem[  1714] = 11'd70;    
		mem[  1715] = 11'd77;    
		mem[  1716] = 11'd35;    
		mem[  1717] = 11'd119;    
		mem[  1718] = 11'd84;    
		mem[  1719] = 11'd40;    
		mem[  1720] = 11'd122;    
		mem[  1721] = 11'd83;    
		mem[  1722] = 11'd41;    
		mem[  1723] = 11'd38;    
		mem[  1724] = 11'd84;    
		mem[  1725] = 11'd83;    
		mem[  1726] = 11'd40;    
		mem[  1727] = 11'd122;    
		mem[  1728] = 11'd41;    
		mem[  1729] = 11'd41;    
		mem[  1730] = 11'd43;    
		mem[  1731] = 11'd40;    
		mem[  1732] = 11'd42;    
		mem[  1733] = 11'd40;    
		mem[  1734] = 11'd42;    
		mem[  1735] = 11'd40;    
		mem[  1736] = 11'd42;    
		mem[  1737] = 11'd39;    
		mem[  1738] = 11'd42;    
		mem[  1739] = 11'd40;    
		mem[  1740] = 11'd42;    
		mem[  1741] = 11'd40;    
		mem[  1742] = 11'd42;    
		mem[  1743] = 11'd35;    
		mem[  1744] = 11'd64;    
		mem[  1745] = 11'd58;    
		mem[  1746] = 11'd54;    
		mem[  1747] = 11'd22;    
		mem[  1748] = 11'd109;    
		mem[  1749] = 11'd59;    
		mem[  1750] = 11'd55;    
		mem[  1751] = 11'd22;    
		mem[  1752] = 11'd109;    
		mem[  1753] = 11'd60;    
		mem[  1754] = 11'd54;    
		mem[  1755] = 11'd22;    
		mem[  1756] = 11'd45;    
		mem[  1757] = 11'd64;    
		mem[  1758] = 11'd60;    
		mem[  1759] = 11'd55;    
		mem[  1760] = 11'd21;    
		mem[  1761] = 11'd45;    
		mem[  1762] = 11'd65;    
		mem[  1763] = 11'd59;    
		mem[  1764] = 11'd58;    
		mem[  1765] = 11'd18;    
		mem[  1766] = 11'd45;    
		mem[  1767] = 11'd64;    
		mem[  1768] = 11'd60;    
		mem[  1769] = 11'd58;    
		mem[  1770] = 11'd18;    
		mem[  1771] = 11'd123;    
		mem[  1772] = 11'd93;    
		mem[  1773] = 11'd32;    
		mem[  1774] = 11'd121;    
		mem[  1775] = 11'd93;    
		mem[  1776] = 11'd32;    
		mem[  1777] = 11'd120;    
		mem[  1778] = 11'd93;    
		mem[  1779] = 11'd31;    
		mem[  1780] = 11'd37;    
		mem[  1781] = 11'd64;    
		mem[  1782] = 11'd28;    
		mem[  1783] = 11'd30;    
		mem[  1784] = 11'd61;    
		mem[  1785] = 11'd31;    
		mem[  1786] = 11'd30;    
		mem[  1787] = 11'd35;    
		mem[  1788] = 11'd29;    
		mem[  1789] = 11'd28;    
		mem[  1790] = 11'd31;    
		mem[  1791] = 11'd35;    
		mem[  1792] = 11'd27;    
		mem[  1793] = 11'd30;    
		mem[  1794] = 11'd18;    
		mem[  1795] = 11'd13;    
		mem[  1796] = 11'd34;    
		mem[  1797] = 11'd29;    
		mem[  1798] = 11'd29;    
		mem[  1799] = 11'd31;    
		mem[  1800] = 11'd35;    
		mem[  1801] = 11'd26;    
		mem[  1802] = 11'd32;    
		mem[  1803] = 11'd30;    
		mem[  1804] = 11'd31;    
		mem[  1805] = 11'd30;    
		mem[  1806] = 11'd31;    
		mem[  1807] = 11'd30;    
		mem[  1808] = 11'd31;    
		mem[  1809] = 11'd31;    
		mem[  1810] = 11'd31;    
		mem[  1811] = 11'd30;    
		mem[  1812] = 11'd31;    
		mem[  1813] = 11'd30;    
		mem[  1814] = 11'd31;    
		mem[  1815] = 11'd30;    
		mem[  1816] = 11'd31;    
		mem[  1817] = 11'd31;    
		mem[  1818] = 11'd31;    
		mem[  1819] = 11'd30;    
		mem[  1820] = 11'd31;    
		mem[  1821] = 11'd30;    
		mem[  1822] = 11'd31;    
		mem[  1823] = 11'd30;    
		mem[  1824] = 11'd32;    
		mem[  1825] = 11'd30;    
		mem[  1826] = 11'd31;    
		mem[  1827] = 11'd30;    
		mem[  1828] = 11'd31;    
		mem[  1829] = 11'd30;    
		mem[  1830] = 11'd32;    
		mem[  1831] = 11'd30;    
		mem[  1832] = 11'd31;    
		mem[  1833] = 11'd30;    
		mem[  1834] = 11'd31;    
		mem[  1835] = 11'd30;    
		mem[  1836] = 11'd31;    
		mem[  1837] = 11'd30;    
		mem[  1838] = 11'd31;    
		mem[  1839] = 11'd31;    
		mem[  1840] = 11'd31;    
		mem[  1841] = 11'd30;    
		mem[  1842] = 11'd31;    
		mem[  1843] = 11'd30;    
		mem[  1844] = 11'd31;    
		mem[  1845] = 11'd31;    
		mem[  1846] = 11'd31;    
		mem[  1847] = 11'd30;    
		mem[  1848] = 11'd31;    
		mem[  1849] = 11'd30;    
		mem[  1850] = 11'd31;    
		mem[  1851] = 11'd30;    
		mem[  1852] = 11'd32;    
		mem[  1853] = 11'd30;    
		mem[  1854] = 11'd31;    
		mem[  1855] = 11'd30;    
		mem[  1856] = 11'd31;    
		mem[  1857] = 11'd30;    
		mem[  1858] = 11'd31;    
		mem[  1859] = 11'd30;    
		mem[  1860] = 11'd32;    
		mem[  1861] = 11'd30;    
		mem[  1862] = 11'd30;    
		mem[  1863] = 11'd31;    
		mem[  1864] = 11'd31;    
		mem[  1865] = 11'd30;    
		mem[  1866] = 11'd31;    
		mem[  1867] = 11'd30;    
		mem[  1868] = 11'd32;    
		mem[  1869] = 11'd30;    
		mem[  1870] = 11'd31;    
		mem[  1871] = 11'd30;    
		mem[  1872] = 11'd31;    
		mem[  1873] = 11'd30;    
		mem[  1874] = 11'd55;    
		mem[  1875] = 11'd57;    
		mem[  1876] = 11'd52;    
		mem[  1877] = 11'd55;    
		mem[  1878] = 11'd29;    
		mem[  1879] = 11'd83;    
		mem[  1880] = 11'd50;    
		mem[  1881] = 11'd59;    
		mem[  1882] = 11'd14;    
		mem[  1883] = 11'd11;    
		mem[  1884] = 11'd28;    
		mem[  1885] = 11'd54;    
		mem[  1886] = 11'd56;    
		mem[  1887] = 11'd52;    
		mem[  1888] = 11'd56;    
		mem[  1889] = 11'd27;    
		mem[  1890] = 11'd79;    
		mem[  1891] = 11'd50;    
		mem[  1892] = 11'd53;    
		mem[  1893] = 11'd27;    
		mem[  1894] = 11'd12;    
		mem[  1895] = 11'd11;    
		mem[  1896] = 11'd12;    
		mem[  1897] = 11'd68;    
		mem[  1898] = 11'd26;    
		mem[  1899] = 11'd25;    
		mem[  1900] = 11'd12;    
		mem[  1901] = 11'd10;    
		mem[  1902] = 11'd56;    
		mem[  1903] = 11'd23;    
		mem[  1904] = 11'd27;    
		mem[  1905] = 11'd50;    
		mem[  1906] = 11'd54;    
		mem[  1907] = 11'd24;    
		mem[  1908] = 11'd79;    
		mem[  1909] = 11'd25;    
		mem[  1910] = 11'd25;    
		mem[  1911] = 11'd26;    
		mem[  1912] = 11'd26;    
		mem[  1913] = 11'd26;    
		mem[  1914] = 11'd26;    
		mem[  1915] = 11'd26;    
		mem[  1916] = 11'd25;    
		mem[  1917] = 11'd26;    
		mem[  1918] = 11'd26;    
		mem[  1919] = 11'd26;    
		mem[  1920] = 11'd25;    
		mem[  1921] = 11'd27;    
		mem[  1922] = 11'd25;    
		mem[  1923] = 11'd26;    
		mem[  1924] = 11'd26;    
		mem[  1925] = 11'd26;    
		mem[  1926] = 11'd25;    
		mem[  1927] = 11'd26;    
		mem[  1928] = 11'd26;    
		mem[  1929] = 11'd26;    
		mem[  1930] = 11'd26;    
		mem[  1931] = 11'd26;    
		mem[  1932] = 11'd25;    
		mem[  1933] = 11'd26;    
		mem[  1934] = 11'd26;    
		mem[  1935] = 11'd26;    
		mem[  1936] = 11'd26;    
		mem[  1937] = 11'd26;    
		mem[  1938] = 11'd24;    
		mem[  1939] = 11'd55;    
		mem[  1940] = 11'd27;    
		mem[  1941] = 11'd20;    
		mem[  1942] = 11'd55;    
		mem[  1943] = 11'd29;    
		mem[  1944] = 11'd10;    
		mem[  1945] = 11'd66;    
		mem[  1946] = 11'd23;    
		mem[  1947] = 11'd77;    
		mem[  1948] = 11'd26;    
		mem[  1949] = 11'd79;    
		mem[  1950] = 11'd50;    
		mem[  1951] = 11'd42;    
		mem[  1952] = 11'd10;    
		mem[  1953] = 11'd50;    
		mem[  1954] = 11'd54;    
		mem[  1955] = 11'd53;    
		mem[  1956] = 11'd24;    
		mem[  1957] = 11'd25;    
		mem[  1958] = 11'd52;    
		mem[  1959] = 11'd51;    
		mem[  1960] = 11'd54;    
		mem[  1961] = 11'd49;    
		mem[  1962] = 11'd54;    
		mem[  1963] = 11'd27;    
		mem[  1964] = 11'd12;    
		mem[  1965] = 11'd9;    
		mem[  1966] = 11'd55;    
		mem[  1967] = 11'd27;    
		mem[  1968] = 11'd21;    
		mem[  1969] = 11'd29;    
		mem[  1970] = 11'd27;    
		mem[  1971] = 11'd24;    
		mem[  1972] = 11'd24;    
		mem[  1973] = 11'd52;    
		mem[  1974] = 11'd26;    
		mem[  1975] = 11'd25;    
		mem[  1976] = 11'd56;    
		mem[  1977] = 11'd47;    
		mem[  1978] = 11'd26;    
		mem[  1979] = 11'd22;    
		mem[  1980] = 11'd26;    
		mem[  1981] = 11'd23;    
		mem[  1982] = 11'd25;    
		mem[  1983] = 11'd24;    
		mem[  1984] = 11'd24;    
		mem[  1985] = 11'd24;    
		mem[  1986] = 11'd25;    
		mem[  1987] = 11'd24;    
		mem[  1988] = 11'd25;    
		mem[  1989] = 11'd24;    
		mem[  1990] = 11'd99;    
		mem[  1991] = 11'd26;    
		mem[  1992] = 11'd74;    
		mem[  1993] = 11'd10;    
		mem[  1994] = 11'd11;    
		mem[  1995] = 11'd73;    
		mem[  1996] = 11'd25;    
		mem[  1997] = 11'd75;    
		mem[  1998] = 11'd44;    
		mem[  1999] = 11'd44;    
		mem[  2000] = 11'd15;    
		mem[  2001] = 11'd33;    
		mem[  2002] = 11'd49;    
		mem[  2003] = 11'd44;    
		mem[  2004] = 11'd44;    
		mem[  2005] = 11'd15;    
		mem[  2006] = 11'd33;    
		mem[  2007] = 11'd49;    
		mem[  2008] = 11'd44;    
		mem[  2009] = 11'd44;    
		mem[  2010] = 11'd15;    
		mem[  2011] = 11'd33;    
		mem[  2012] = 11'd49;    
		mem[  2013] = 11'd44;    
		mem[  2014] = 11'd44;    
		mem[  2015] = 11'd15;    
		mem[  2016] = 11'd33;    
		mem[  2017] = 11'd49;    
		mem[  2018] = 11'd44;    
		mem[  2019] = 11'd44;    
		mem[  2020] = 11'd14;    
		mem[  2021] = 11'd34;    
		mem[  2022] = 11'd49;    
		mem[  2023] = 11'd44;    
		mem[  2024] = 11'd44;    
		mem[  2025] = 11'd14;    
		mem[  2026] = 11'd34;    
		mem[  2027] = 11'd48;    
		mem[  2028] = 11'd24;    
		mem[  2029] = 11'd22;    
		mem[  2030] = 11'd24;    
		mem[  2031] = 11'd22;    
		mem[  2032] = 11'd23;    
		mem[  2033] = 11'd23;    
		mem[  2034] = 11'd23;    
		mem[  2035] = 11'd23;    
		mem[  2036] = 11'd23;    
		mem[  2037] = 11'd23;    
		mem[  2038] = 11'd23;    
		mem[  2039] = 11'd23;    
		mem[  2040] = 11'd24;    
		mem[  2041] = 11'd23;    
		mem[  2042] = 11'd25;    
		mem[  2043] = 11'd21;    
		mem[  2044] = 11'd47;    
		mem[  2045] = 11'd23;    
		mem[  2046] = 11'd22;    
		mem[  2047] = 11'd47;    
		mem[  2048] = 11'd45;    
		mem[  2049] = 11'd49;    
		mem[  2050] = 11'd43;    
		mem[  2051] = 11'd50;    
		mem[  2052] = 11'd23;    
		mem[  2053] = 11'd11;    
		mem[  2054] = 11'd57;    
		mem[  2055] = 11'd24;    
		mem[  2056] = 11'd46;    
		mem[  2057] = 11'd24;    
		mem[  2058] = 11'd21;    
		mem[  2059] = 11'd21;    
		mem[  2060] = 11'd46;    
		mem[  2061] = 11'd15;    
		mem[  2062] = 11'd32;    
		mem[  2063] = 11'd49;    
		mem[  2064] = 11'd46;    
		mem[  2065] = 11'd24;    
		mem[  2066] = 11'd22;    
		mem[  2067] = 11'd45;    
		mem[  2068] = 11'd46;    
		mem[  2069] = 11'd49;    
		mem[  2070] = 11'd9;    
		mem[  2071] = 11'd10;    
		mem[  2072] = 11'd24;    
		mem[  2073] = 11'd49;    
		mem[  2074] = 11'd43;    
		mem[  2075] = 11'd49;    
		mem[  2076] = 11'd26;    
		mem[  2077] = 11'd9;    
		mem[  2078] = 11'd8;    
		mem[  2079] = 11'd50;    
		mem[  2080] = 11'd21;    
		mem[  2081] = 11'd69;    
		mem[  2082] = 11'd23;    
		mem[  2083] = 11'd71;    
		mem[  2084] = 11'd443;    
		mem[  2085] = 11'd21;    
		mem[  2086] = 11'd80;    
		mem[  2087] = 11'd60;    
		mem[  2088] = 11'd20;    
		mem[  2089] = 11'd80;    
		mem[  2090] = 11'd67;    
		mem[  2091] = 11'd95;    
		mem[  2092] = 11'd48;    
		mem[  2093] = 11'd20;    
		mem[  2094] = 11'd24;    
		mem[  2095] = 11'd49;    
		mem[  2096] = 11'd23;    
		mem[  2097] = 11'd67;    
		mem[  2098] = 11'd22;    
		mem[  2099] = 11'd72;    
		mem[  2100] = 11'd47;    
		mem[  2101] = 11'd21;    
		mem[  2102] = 11'd23;    
		mem[  2103] = 11'd48;    
		mem[  2104] = 11'd24;    
		mem[  2105] = 11'd11;    
		mem[  2106] = 11'd56;    
		mem[  2107] = 11'd23;    
		mem[  2108] = 11'd70;    
		mem[  2109] = 11'd42;    
		mem[  2110] = 11'd24;    
		mem[  2111] = 11'd10;    
		mem[  2112] = 11'd10;    
		mem[  2113] = 11'd43;    
		mem[  2114] = 11'd44;    
		mem[  2115] = 11'd45;    
		mem[  2116] = 11'd20;    
		mem[  2117] = 11'd22;    
		mem[  2118] = 11'd44;    
		mem[  2119] = 11'd42;    
		mem[  2120] = 11'd44;    
		mem[  2121] = 11'd43;    
		mem[  2122] = 11'd22;    
		mem[  2123] = 11'd22;    
		mem[  2124] = 11'd22;    
		mem[  2125] = 11'd22;    
		mem[  2126] = 11'd22;    
		mem[  2127] = 11'd22;    
		mem[  2128] = 11'd22;    
		mem[  2129] = 11'd21;    
		mem[  2130] = 11'd23;    
		mem[  2131] = 11'd21;    
		mem[  2132] = 11'd22;    
		mem[  2133] = 11'd22;    
		mem[  2134] = 11'd54;    
		mem[  2135] = 11'd31;    
		mem[  2136] = 11'd45;    
		mem[  2137] = 11'd44;    
		mem[  2138] = 11'd21;    
		mem[  2139] = 11'd21;    
		mem[  2140] = 11'd43;    
		mem[  2141] = 11'd43;    
		mem[  2142] = 11'd47;    
		mem[  2143] = 11'd23;    
		mem[  2144] = 11'd52;    
		mem[  2145] = 11'd12;    
		mem[  2146] = 11'd44;    
		mem[  2147] = 11'd20;    
		mem[  2148] = 11'd22;    
		mem[  2149] = 11'd22;    
		mem[  2150] = 11'd21;    
		mem[  2151] = 11'd46;    
		mem[  2152] = 11'd44;    
		mem[  2153] = 11'd32;    
		mem[  2154] = 11'd53;    
		mem[  2155] = 11'd45;    
		mem[  2156] = 11'd20;    
		mem[  2157] = 11'd65;    
		mem[  2158] = 11'd44;    
		mem[  2159] = 11'd11;    
		mem[  2160] = 11'd33;    
		mem[  2161] = 11'd34;    
		mem[  2162] = 11'd45;    
		mem[  2163] = 11'd10;    
		mem[  2164] = 11'd43;    
		mem[  2165] = 11'd21;    
		mem[  2166] = 11'd20;    
		mem[  2167] = 11'd24;    
		mem[  2168] = 11'd20;    
		mem[  2169] = 11'd46;    
		mem[  2170] = 11'd43;    
		mem[  2171] = 11'd18;    
		mem[  2172] = 11'd23;    
		mem[  2173] = 11'd46;    
		mem[  2174] = 11'd44;    
		mem[  2175] = 11'd21;    
		mem[  2176] = 11'd64;    
		mem[  2177] = 11'd23;    
		mem[  2178] = 11'd21;    
		mem[  2179] = 11'd20;    
		mem[  2180] = 11'd23;    
		mem[  2181] = 11'd43;    
		mem[  2182] = 11'd44;    
		mem[  2183] = 11'd45;    
		mem[  2184] = 11'd22;    
		mem[  2185] = 11'd20;    
		mem[  2186] = 11'd25;    
		mem[  2187] = 11'd20;    
		mem[  2188] = 11'd45;    
		mem[  2189] = 11'd19;    
		mem[  2190] = 11'd23;    
		mem[  2191] = 11'd21;    
		mem[  2192] = 11'd21;    
		mem[  2193] = 11'd23;    
		mem[  2194] = 11'd23;    
		mem[  2195] = 11'd44;    
		mem[  2196] = 11'd23;    
		mem[  2197] = 11'd9;    
		mem[  2198] = 11'd8;    
		mem[  2199] = 11'd45;    
		mem[  2200] = 11'd45;    
		mem[  2201] = 11'd20;    
		mem[  2202] = 11'd22;    
		mem[  2203] = 11'd43;    
		mem[  2204] = 11'd43;    
		mem[  2205] = 11'd46;    
		mem[  2206] = 11'd23;    
		mem[  2207] = 11'd10;    
		mem[  2208] = 11'd8;    
		mem[  2209] = 11'd35;    
		mem[  2210] = 11'd11;    
		mem[  2211] = 11'd44;    
		mem[  2212] = 11'd20;    
		mem[  2213] = 11'd22;    
		mem[  2214] = 11'd23;    
		mem[  2215] = 11'd20;    
		mem[  2216] = 11'd45;    
		mem[  2217] = 11'd44;    
		mem[  2218] = 11'd42;    
		mem[  2219] = 11'd24;    
		mem[  2220] = 11'd21;    
		mem[  2221] = 11'd44;    
		mem[  2222] = 11'd21;    
		mem[  2223] = 11'd21;    
		mem[  2224] = 11'd43;    
		mem[  2225] = 11'd25;    
		mem[  2226] = 11'd19;    
		mem[  2227] = 11'd21;    
		mem[  2228] = 11'd23;    
		mem[  2229] = 11'd35;    
		mem[  2230] = 11'd45;    
		mem[  2231] = 11'd9;    
		mem[  2232] = 11'd43;    
		mem[  2233] = 11'd21;    
		mem[  2234] = 11'd20;    
		mem[  2235] = 11'd25;    
		mem[  2236] = 11'd19;    
		mem[  2237] = 11'd47;    
		mem[  2238] = 11'd43;    
		mem[  2239] = 11'd17;    
		mem[  2240] = 11'd22;    
		mem[  2241] = 11'd47;    
		mem[  2242] = 11'd44;    
		mem[  2243] = 11'd22;    
		mem[  2244] = 11'd63;    
		mem[  2245] = 11'd44;    
		mem[  2246] = 11'd20;    
		mem[  2247] = 11'd23;    
		mem[  2248] = 11'd42;    
		mem[  2249] = 11'd45;    
		mem[  2250] = 11'd46;    
		mem[  2251] = 11'd27;    
		mem[  2252] = 11'd11;    
		mem[  2253] = 11'd59;    
		mem[  2254] = 11'd23;    
		mem[  2255] = 11'd75;    
		mem[  2256] = 11'd51;    
		mem[  2257] = 11'd44;    
		mem[  2258] = 11'd54;    
		mem[  2259] = 11'd21;    
		mem[  2260] = 11'd25;    
		mem[  2261] = 11'd37;    
		mem[  2262] = 11'd14;    
		mem[  2263] = 11'd48;    
		mem[  2264] = 11'd46;    
		mem[  2265] = 11'd51;    
		mem[  2266] = 11'd24;    
		mem[  2267] = 11'd75;    
		mem[  2268] = 11'd49;    
		mem[  2269] = 11'd20;    
		mem[  2270] = 11'd24;    
		mem[  2271] = 11'd49;    
		mem[  2272] = 11'd23;    
		mem[  2273] = 11'd67;    
		mem[  2274] = 11'd22;    
		mem[  2275] = 11'd23;    
		mem[  2276] = 11'd49;    
		mem[  2277] = 11'd47;    
		mem[  2278] = 11'd21;    
		mem[  2279] = 11'd23;    
		mem[  2280] = 11'd48;    
		mem[  2281] = 11'd24;    
		mem[  2282] = 11'd11;    
		mem[  2283] = 11'd8;    
		mem[  2284] = 11'd48;    
		mem[  2285] = 11'd23;    
		mem[  2286] = 11'd71;    
		mem[  2287] = 11'd46;    
		mem[  2288] = 11'd23;    
		mem[  2289] = 11'd22;    
		mem[  2290] = 11'd45;    
		mem[  2291] = 11'd47;    
		mem[  2292] = 11'd23;    
		mem[  2293] = 11'd23;    
		mem[  2294] = 11'd23;    
		mem[  2295] = 11'd24;    
		mem[  2296] = 11'd23;    
		mem[  2297] = 11'd23;    
		mem[  2298] = 11'd24;    
		mem[  2299] = 11'd22;    
		mem[  2300] = 11'd24;    
		mem[  2301] = 11'd23;    
		mem[  2302] = 11'd23;    
		mem[  2303] = 11'd23;    
		mem[  2304] = 11'd24;    
		mem[  2305] = 11'd67;    
		mem[  2306] = 11'd49;    
		mem[  2307] = 11'd35;    
		mem[  2308] = 11'd8;    
		mem[  2309] = 11'd51;    
		mem[  2310] = 11'd20;    
		mem[  2311] = 11'd69;    
		mem[  2312] = 11'd22;    
		mem[  2313] = 11'd72;    
		mem[  2314] = 11'd45;    
		mem[  2315] = 11'd26;    
		mem[  2316] = 11'd9;    
		mem[  2317] = 11'd12;    
		mem[  2318] = 11'd45;    
		mem[  2319] = 11'd47;    
		mem[  2320] = 11'd48;    
		mem[  2321] = 11'd21;    
		mem[  2322] = 11'd23;    
		mem[  2323] = 11'd47;    
		mem[  2324] = 11'd44;    
		mem[  2325] = 11'd49;    
		mem[  2326] = 11'd36;    
		mem[  2327] = 11'd8;    
		mem[  2328] = 11'd49;    
		mem[  2329] = 11'd23;    
		mem[  2330] = 11'd68;    
		mem[  2331] = 11'd23;    
		mem[  2332] = 11'd71;    
		mem[  2333] = 11'd19;    
		mem[  2334] = 11'd25;    
		mem[  2335] = 11'd46;    
		mem[  2336] = 11'd46;    
		mem[  2337] = 11'd48;    
		mem[  2338] = 11'd47;    
		mem[  2339] = 11'd22;    
		mem[  2340] = 11'd23;    
		mem[  2341] = 11'd46;    
		mem[  2342] = 11'd46;    
		mem[  2343] = 11'd23;    
		mem[  2344] = 11'd23;    
		mem[  2345] = 11'd24;    
		mem[  2346] = 11'd23;    
		mem[  2347] = 11'd23;    
		mem[  2348] = 11'd23;    
		mem[  2349] = 11'd23;    
		mem[  2350] = 11'd23;    
		mem[  2351] = 11'd23;    
		mem[  2352] = 11'd23;    
		mem[  2353] = 11'd24;    
		mem[  2354] = 11'd23;    
		mem[  2355] = 11'd23;    
		mem[  2356] = 11'd23;    
		mem[  2357] = 11'd23;    
		mem[  2358] = 11'd22;    
		mem[  2359] = 11'd58;    
		mem[  2360] = 11'd27;    
		mem[  2361] = 11'd82;    
		mem[  2362] = 11'd56;    
		mem[  2363] = 11'd24;    
		mem[  2364] = 11'd27;    
		mem[  2365] = 11'd59;    
		mem[  2366] = 11'd25;    
		mem[  2367] = 11'd78;    
		mem[  2368] = 11'd15;    
		mem[  2369] = 11'd42;    
		mem[  2370] = 11'd55;    
		mem[  2371] = 11'd57;    
		mem[  2372] = 11'd31;    
		mem[  2373] = 11'd10;    
		mem[  2374] = 11'd40;    
		mem[  2375] = 11'd28;    
		mem[  2376] = 11'd51;    
		mem[  2377] = 11'd29;    
		mem[  2378] = 11'd10;    
		mem[  2379] = 11'd14;    
		mem[  2380] = 11'd50;    
		mem[  2381] = 11'd51;    
		mem[  2382] = 11'd54;    
		mem[  2383] = 11'd48;    
		mem[  2384] = 11'd56;    
		mem[  2385] = 11'd10;    
		mem[  2386] = 11'd13;    
		mem[  2387] = 11'd24;    
		mem[  2388] = 11'd51;    
		mem[  2389] = 11'd15;    
		mem[  2390] = 11'd38;    
		mem[  2391] = 11'd53;    
		mem[  2392] = 11'd53;    
		mem[  2393] = 11'd12;    
		mem[  2394] = 11'd11;    
		mem[  2395] = 11'd26;    
		mem[  2396] = 11'd54;    
		mem[  2397] = 11'd52;    
		mem[  2398] = 11'd51;    
		mem[  2399] = 11'd26;    
		mem[  2400] = 11'd25;    
		mem[  2401] = 11'd26;    
		mem[  2402] = 11'd25;    
		mem[  2403] = 11'd26;    
		mem[  2404] = 11'd25;    
		mem[  2405] = 11'd26;    
		mem[  2406] = 11'd26;    
		mem[  2407] = 11'd26;    
		mem[  2408] = 11'd25;    
		mem[  2409] = 11'd105;    
		mem[  2410] = 11'd48;    
		mem[  2411] = 11'd56;    
		mem[  2412] = 11'd48;    
		mem[  2413] = 11'd56;    
		mem[  2414] = 11'd48;    
		mem[  2415] = 11'd55;    
		mem[  2416] = 11'd48;    
		mem[  2417] = 11'd55;    
		mem[  2418] = 11'd48;    
		mem[  2419] = 11'd55;    
		mem[  2420] = 11'd48;    
		mem[  2421] = 11'd55;    
		mem[  2422] = 11'd49;    
		mem[  2423] = 11'd55;    
		mem[  2424] = 11'd48;    
		mem[  2425] = 11'd55;    
		mem[  2426] = 11'd48;    
		mem[  2427] = 11'd55;    
		mem[  2428] = 11'd48;    
		mem[  2429] = 11'd55;    
		mem[  2430] = 11'd49;    
		mem[  2431] = 11'd54;    
		mem[  2432] = 11'd49;    
		mem[  2433] = 11'd54;    
		mem[  2434] = 11'd49;    
		mem[  2435] = 11'd55;    
		mem[  2436] = 11'd51;    
		mem[  2437] = 11'd27;    
		mem[  2438] = 11'd24;    
		mem[  2439] = 11'd26;    
		mem[  2440] = 11'd25;    
		mem[  2441] = 11'd26;    
		mem[  2442] = 11'd25;    
		mem[  2443] = 11'd26;    
		mem[  2444] = 11'd26;    
		mem[  2445] = 11'd26;    
		mem[  2446] = 11'd26;    
		mem[  2447] = 11'd25;    
		mem[  2448] = 11'd26;    
		mem[  2449] = 11'd26;    
		mem[  2450] = 11'd92;    
		mem[  2451] = 11'd58;    
		mem[  2452] = 11'd64;    
		mem[  2453] = 11'd58;    
		mem[  2454] = 11'd66;    
		mem[  2455] = 11'd57;    
		mem[  2456] = 11'd65;    
		mem[  2457] = 11'd58;    
		mem[  2458] = 11'd65;    
		mem[  2459] = 11'd58;    
		mem[  2460] = 11'd64;    
		mem[  2461] = 11'd58;    
		mem[  2462] = 11'd65;    
		mem[  2463] = 11'd58;    
		mem[  2464] = 11'd64;    
		mem[  2465] = 11'd58;    
		mem[  2466] = 11'd65;    
		mem[  2467] = 11'd58;    
		mem[  2468] = 11'd64;    
		mem[  2469] = 11'd58;    
		mem[  2470] = 11'd65;    
		mem[  2471] = 11'd58;    
		mem[  2472] = 11'd64;    
		mem[  2473] = 11'd61;    
		mem[  2474] = 11'd32;    
		mem[  2475] = 11'd28;    
		mem[  2476] = 11'd32;    
		mem[  2477] = 11'd29;    
		mem[  2478] = 11'd31;    
		mem[  2479] = 11'd30;    
		mem[  2480] = 11'd31;    
		mem[  2481] = 11'd30;    
		mem[  2482] = 11'd31;    
		mem[  2483] = 11'd31;    
		mem[  2484] = 11'd30;    
		mem[  2485] = 11'd94;    
		mem[  2486] = 11'd59;    
		mem[  2487] = 11'd63;    
		mem[  2488] = 11'd60;    
		mem[  2489] = 11'd64;    
		mem[  2490] = 11'd32;    
		mem[  2491] = 11'd10;    
		mem[  2492] = 11'd19;    
		mem[  2493] = 11'd58;    
		mem[  2494] = 11'd64;    
		mem[  2495] = 11'd59;    
		mem[  2496] = 11'd60;    
		mem[  2497] = 11'd32;    
		mem[  2498] = 11'd64;    
		mem[  2499] = 11'd31;    
		mem[  2500] = 11'd13;    
		mem[  2501] = 11'd15;    
		mem[  2502] = 11'd93;    
		mem[  2503] = 11'd36;    
		mem[  2504] = 11'd11;    
		mem[  2505] = 11'd11;    
		mem[  2506] = 11'd66;    
		mem[  2507] = 11'd33;    
		mem[  2508] = 11'd24;    
		mem[  2509] = 11'd65;    
		mem[  2510] = 11'd25;    
		mem[  2511] = 11'd34;    
		mem[  2512] = 11'd62;    
		mem[  2513] = 11'd61;    
		mem[  2514] = 11'd63;    
		mem[  2515] = 11'd31;    
		mem[  2516] = 11'd30;    
		mem[  2517] = 11'd29;    
		mem[  2518] = 11'd31;    
		mem[  2519] = 11'd30;    
		mem[  2520] = 11'd31;    
		mem[  2521] = 11'd31;    
		mem[  2522] = 11'd30;    
		mem[  2523] = 11'd31;    
		mem[  2524] = 11'd30;    
		mem[  2525] = 11'd31;    
		mem[  2526] = 11'd31;    
		mem[  2527] = 11'd31;    
		mem[  2528] = 11'd30;    
		mem[  2529] = 11'd54;    
		mem[  2530] = 11'd59;    
		mem[  2531] = 11'd26;    
		mem[  2532] = 11'd83;    
		mem[  2533] = 11'd24;    
		mem[  2534] = 11'd30;    
		mem[  2535] = 11'd51;    
		mem[  2536] = 11'd59;    
		mem[  2537] = 11'd26;    
		mem[  2538] = 11'd14;    
		mem[  2539] = 11'd9;    
		mem[  2540] = 11'd60;    
		mem[  2541] = 11'd26;    
		mem[  2542] = 11'd28;    
		mem[  2543] = 11'd82;    
		mem[  2544] = 11'd28;    
		mem[  2545] = 11'd26;    
		mem[  2546] = 11'd24;    
		mem[  2547] = 11'd57;    
		mem[  2548] = 11'd26;    
		mem[  2549] = 11'd13;    
		mem[  2550] = 11'd26;    
		mem[  2551] = 11'd9;    
		mem[  2552] = 11'd25;    
		mem[  2553] = 11'd56;    
		mem[  2554] = 11'd49;    
		mem[  2555] = 11'd52;    
		mem[  2556] = 11'd52;    
		mem[  2557] = 11'd50;    
		mem[  2558] = 11'd53;    
		mem[  2559] = 11'd53;    
		mem[  2560] = 11'd24;    
		mem[  2561] = 11'd79;    
		mem[  2562] = 11'd24;    
		mem[  2563] = 11'd27;    
		mem[  2564] = 11'd50;    
		mem[  2565] = 11'd54;    
		mem[  2566] = 11'd26;    
		mem[  2567] = 11'd23;    
		mem[  2568] = 11'd54;    
		mem[  2569] = 11'd27;    
		mem[  2570] = 11'd21;    
		mem[  2571] = 11'd28;    
		mem[  2572] = 11'd24;    
		mem[  2573] = 11'd55;    
		mem[  2574] = 11'd51;    
		mem[  2575] = 11'd50;    
		mem[  2576] = 11'd53;    
		mem[  2577] = 11'd25;    
		mem[  2578] = 11'd25;    
		mem[  2579] = 11'd52;    
		mem[  2580] = 11'd54;    
		mem[  2581] = 11'd24;    
		mem[  2582] = 11'd24;    
		mem[  2583] = 11'd29;    
		mem[  2584] = 11'd26;    
		mem[  2585] = 11'd24;    
		mem[  2586] = 11'd27;    
		mem[  2587] = 11'd50;    
		mem[  2588] = 11'd28;    
		mem[  2589] = 11'd26;    
		mem[  2590] = 11'd26;    
		mem[  2591] = 11'd23;    
		mem[  2592] = 11'd54;    
		mem[  2593] = 11'd28;    
		mem[  2594] = 11'd21;    
		mem[  2595] = 11'd27;    
		mem[  2596] = 11'd15;    
		mem[  2597] = 11'd10;    
		mem[  2598] = 11'd53;    
		mem[  2599] = 11'd52;    
		mem[  2600] = 11'd50;    
		mem[  2601] = 11'd30;    
		mem[  2602] = 11'd23;    
		mem[  2603] = 11'd51;    
		mem[  2604] = 11'd51;    
		mem[  2605] = 11'd30;    
		mem[  2606] = 11'd23;    
		mem[  2607] = 11'd25;    
		mem[  2608] = 11'd25;    
		mem[  2609] = 11'd25;    
		mem[  2610] = 11'd27;    
		mem[  2611] = 11'd26;    
		mem[  2612] = 11'd26;    
		mem[  2613] = 11'd26;    
		mem[  2614] = 11'd26;    
		mem[  2615] = 11'd26;    
		mem[  2616] = 11'd25;    
		mem[  2617] = 11'd26;    
		mem[  2618] = 11'd26;    
		mem[  2619] = 11'd26;    
		mem[  2620] = 11'd26;    
		mem[  2621] = 11'd26;    
		mem[  2622] = 11'd25;    
		mem[  2623] = 11'd27;    
		mem[  2624] = 11'd25;    
		mem[  2625] = 11'd26;    
		mem[  2626] = 11'd25;    
		mem[  2627] = 11'd27;    
		mem[  2628] = 11'd25;    
		mem[  2629] = 11'd26;    
		mem[  2630] = 11'd26;    
		mem[  2631] = 11'd26;    
		mem[  2632] = 11'd25;    
		mem[  2633] = 11'd26;    
		mem[  2634] = 11'd26;    
		mem[  2635] = 11'd26;    
		mem[  2636] = 11'd25;    
		mem[  2637] = 11'd27;    
		mem[  2638] = 11'd52;    
		mem[  2639] = 11'd27;    
		mem[  2640] = 11'd48;    
		mem[  2641] = 11'd56;    
		mem[  2642] = 11'd24;    
		mem[  2643] = 11'd15;    
		mem[  2644] = 11'd7;    
		mem[  2645] = 11'd56;    
		mem[  2646] = 11'd25;    
		mem[  2647] = 11'd25;    
		mem[  2648] = 11'd78;    
		mem[  2649] = 11'd27;    
		mem[  2650] = 11'd26;    
		mem[  2651] = 11'd22;    
		mem[  2652] = 11'd55;    
		mem[  2653] = 11'd26;    
		mem[  2654] = 11'd10;    
		mem[  2655] = 11'd14;    
		mem[  2656] = 11'd79;    
		mem[  2657] = 11'd26;    
		mem[  2658] = 11'd27;    
		mem[  2659] = 11'd21;    
		mem[  2660] = 11'd55;    
		mem[  2661] = 11'd26;    
		mem[  2662] = 11'd12;    
		mem[  2663] = 11'd12;    
		mem[  2664] = 11'd12;    
		mem[  2665] = 11'd66;    
		mem[  2666] = 11'd27;    
		mem[  2667] = 11'd28;    
		mem[  2668] = 11'd20;    
		mem[  2669] = 11'd55;    
		mem[  2670] = 11'd27;    
		mem[  2671] = 11'd13;    
		mem[  2672] = 11'd34;    
		mem[  2673] = 11'd25;    
		mem[  2674] = 11'd28;    
		mem[  2675] = 11'd28;    
		mem[  2676] = 11'd49;    
		mem[  2677] = 11'd54;    
		mem[  2678] = 11'd27;    
		mem[  2679] = 11'd15;    
		mem[  2680] = 11'd33;    
		mem[  2681] = 11'd25;    
		mem[  2682] = 11'd34;    
		mem[  2683] = 11'd33;    
		mem[  2684] = 11'd30;    
		mem[  2685] = 11'd30;    
		mem[  2686] = 11'd67;    
		mem[  2687] = 11'd34;    
		mem[  2688] = 11'd29;    
		mem[  2689] = 11'd36;    
		mem[  2690] = 11'd34;    
		mem[  2691] = 11'd30;    
		mem[  2692] = 11'd30;    
		mem[  2693] = 11'd67;    
		mem[  2694] = 11'd33;    
		mem[  2695] = 11'd30;    
		mem[  2696] = 11'd36;    
		mem[  2697] = 11'd33;    
		mem[  2698] = 11'd31;    
		mem[  2699] = 11'd30;    
		mem[  2700] = 11'd67;    
		mem[  2701] = 11'd33;    
		mem[  2702] = 11'd16;    
		mem[  2703] = 11'd12;    
		mem[  2704] = 11'd32;    
		mem[  2705] = 11'd33;    
		mem[  2706] = 11'd30;    
		mem[  2707] = 11'd17;    
		mem[  2708] = 11'd11;    
		mem[  2709] = 11'd34;    
		mem[  2710] = 11'd30;    
		mem[  2711] = 11'd59;    
		mem[  2712] = 11'd63;    
		mem[  2713] = 11'd32;    
		mem[  2714] = 11'd28;    
		mem[  2715] = 11'd63;    
		mem[  2716] = 11'd29;    
		mem[  2717] = 11'd31;    
		mem[  2718] = 11'd61;    
		mem[  2719] = 11'd34;    
		mem[  2720] = 11'd28;    
		mem[  2721] = 11'd61;    
		mem[  2722] = 11'd62;    
		mem[  2723] = 11'd33;    
		mem[  2724] = 11'd28;    
		mem[  2725] = 11'd31;    
		mem[  2726] = 11'd30;    
		mem[  2727] = 11'd31;    
		mem[  2728] = 11'd30;    
		mem[  2729] = 11'd30;    
		mem[  2730] = 11'd31;    
		mem[  2731] = 11'd30;    
		mem[  2732] = 11'd31;    
		mem[  2733] = 11'd30;    
		mem[  2734] = 11'd31;    
		mem[  2735] = 11'd31;    
		mem[  2736] = 11'd30;    
		mem[  2737] = 11'd31;    
		mem[  2738] = 11'd31;    
		mem[  2739] = 11'd31;    
		mem[  2740] = 11'd30;    
		mem[  2741] = 11'd31;    
		mem[  2742] = 11'd30;    
		mem[  2743] = 11'd31;    
		mem[  2744] = 11'd31;    
		mem[  2745] = 11'd29;    
		mem[  2746] = 11'd33;    
		mem[  2747] = 11'd59;    
		mem[  2748] = 11'd63;    
		mem[  2749] = 11'd63;    
		mem[  2750] = 11'd31;    
		mem[  2751] = 11'd30;    
		mem[  2752] = 11'd59;    
		mem[  2753] = 11'd63;    
		mem[  2754] = 11'd62;    
		mem[  2755] = 11'd31;    
		mem[  2756] = 11'd30;    
		mem[  2757] = 11'd59;    
		mem[  2758] = 11'd62;    
		mem[  2759] = 11'd63;    
		mem[  2760] = 11'd31;    
		mem[  2761] = 11'd30;    
		mem[  2762] = 11'd59;    
		mem[  2763] = 11'd63;    
		mem[  2764] = 11'd62;    
		mem[  2765] = 11'd31;    
		mem[  2766] = 11'd30;    
		mem[  2767] = 11'd59;    
		mem[  2768] = 11'd63;    
		mem[  2769] = 11'd62;    
		mem[  2770] = 11'd31;    
		mem[  2771] = 11'd30;    
		mem[  2772] = 11'd60;    
		mem[  2773] = 11'd62;    
		mem[  2774] = 11'd62;    
		mem[  2775] = 11'd31;    
		mem[  2776] = 11'd30;    
		mem[  2777] = 11'd59;    
		mem[  2778] = 11'd63;    
		mem[  2779] = 11'd62;    
		mem[  2780] = 11'd31;    
		mem[  2781] = 11'd30;    
		mem[  2782] = 11'd60;    
		mem[  2783] = 11'd62;    
		mem[  2784] = 11'd62;    
		mem[  2785] = 11'd31;    
		mem[  2786] = 11'd30;    
		mem[  2787] = 11'd60;    
		mem[  2788] = 11'd62;    
		mem[  2789] = 11'd62;    
		mem[  2790] = 11'd31;    
		mem[  2791] = 11'd30;    
		mem[  2792] = 11'd60;    
		mem[  2793] = 11'd62;    
		mem[  2794] = 11'd62;    
		mem[  2795] = 11'd31;    
		mem[  2796] = 11'd30;    
		mem[  2797] = 11'd60;    
		mem[  2798] = 11'd62;    
		mem[  2799] = 11'd62;    
		mem[  2800] = 11'd31;    
		mem[  2801] = 11'd30;    
		mem[  2802] = 11'd60;    
		mem[  2803] = 11'd62;    
		mem[  2804] = 11'd63;    
		mem[  2805] = 11'd31;    
		mem[  2806] = 11'd30;    
		mem[  2807] = 11'd59;    
		mem[  2808] = 11'd62;    
		mem[  2809] = 11'd63;    
		mem[  2810] = 11'd31;    
		mem[  2811] = 11'd30;    
		mem[  2812] = 11'd59;    
		mem[  2813] = 11'd62;    
		mem[  2814] = 11'd63;    
		mem[  2815] = 11'd31;    
		mem[  2816] = 11'd30;    
		mem[  2817] = 11'd59;    
		mem[  2818] = 11'd62;    
		mem[  2819] = 11'd63;    
		mem[  2820] = 11'd31;    
		mem[  2821] = 11'd30;    
		mem[  2822] = 11'd59;    
		mem[  2823] = 11'd62;    
		mem[  2824] = 11'd63;    
		mem[  2825] = 11'd31;    
		mem[  2826] = 11'd30;    
		mem[  2827] = 11'd59;    
		mem[  2828] = 11'd62;    
		mem[  2829] = 11'd63;    
		mem[  2830] = 11'd31;    
		mem[  2831] = 11'd30;    
		mem[  2832] = 11'd59;    
		mem[  2833] = 11'd62;    

	end
	
endmodule
