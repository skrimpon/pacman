module pacman_extrapac_converted(in, out, clk); //ok
	 input [10:0] in;
	 input clk;
	 output reg [6:0] out;
	 
	 reg  [6:0] mem [0:1394];
	 always @(posedge clk) out  =  mem[ in ];
	 
	 initial begin
		mem[     0] = 7'd26;    
		mem[     1] = 7'd44;    
		mem[     2] = 7'd13;    
		mem[     3] = 7'd17;    
		mem[     4] = 7'd28;    
		mem[     5] = 7'd29;    
		mem[     6] = 7'd29;    
		mem[     7] = 7'd30;    
		mem[     8] = 7'd29;    
		mem[     9] = 7'd30;    
		mem[    10] = 7'd29;    
		mem[    11] = 7'd29;    
		mem[    12] = 7'd30;    
		mem[    13] = 7'd29;    
		mem[    14] = 7'd30;    
		mem[    15] = 7'd29;    
		mem[    16] = 7'd29;    
		mem[    17] = 7'd30;    
		mem[    18] = 7'd29;    
		mem[    19] = 7'd30;    
		mem[    20] = 7'd29;    
		mem[    21] = 7'd30;    
		mem[    22] = 7'd29;    
		mem[    23] = 7'd30;    
		mem[    24] = 7'd29;    
		mem[    25] = 7'd29;    
		mem[    26] = 7'd30;    
		mem[    27] = 7'd29;    
		mem[    28] = 7'd30;    
		mem[    29] = 7'd29;    
		mem[    30] = 7'd30;    
		mem[    31] = 7'd29;    
		mem[    32] = 7'd30;    
		mem[    33] = 7'd29;    
		mem[    34] = 7'd30;    
		mem[    35] = 7'd29;    
		mem[    36] = 7'd29;    
		mem[    37] = 7'd30;    
		mem[    38] = 7'd29;    
		mem[    39] = 7'd30;    
		mem[    40] = 7'd29;    
		mem[    41] = 7'd30;    
		mem[    42] = 7'd29;    
		mem[    43] = 7'd30;    
		mem[    44] = 7'd29;    
		mem[    45] = 7'd30;    
		mem[    46] = 7'd29;    
		mem[    47] = 7'd29;    
		mem[    48] = 7'd30;    
		mem[    49] = 7'd29;    
		mem[    50] = 7'd30;    
		mem[    51] = 7'd29;    
		mem[    52] = 7'd30;    
		mem[    53] = 7'd29;    
		mem[    54] = 7'd29;    
		mem[    55] = 7'd30;    
		mem[    56] = 7'd29;    
		mem[    57] = 7'd30;    
		mem[    58] = 7'd29;    
		mem[    59] = 7'd30;    
		mem[    60] = 7'd29;    
		mem[    61] = 7'd30;    
		mem[    62] = 7'd29;    
		mem[    63] = 7'd29;    
		mem[    64] = 7'd30;    
		mem[    65] = 7'd29;    
		mem[    66] = 7'd30;    
		mem[    67] = 7'd29;    
		mem[    68] = 7'd30;    
		mem[    69] = 7'd29;    
		mem[    70] = 7'd30;    
		mem[    71] = 7'd29;    
		mem[    72] = 7'd29;    
		mem[    73] = 7'd30;    
		mem[    74] = 7'd29;    
		mem[    75] = 7'd30;    
		mem[    76] = 7'd29;    
		mem[    77] = 7'd30;    
		mem[    78] = 7'd29;    
		mem[    79] = 7'd30;    
		mem[    80] = 7'd29;    
		mem[    81] = 7'd30;    
		mem[    82] = 7'd29;    
		mem[    83] = 7'd29;    
		mem[    84] = 7'd30;    
		mem[    85] = 7'd29;    
		mem[    86] = 7'd30;    
		mem[    87] = 7'd29;    
		mem[    88] = 7'd29;    
		mem[    89] = 7'd30;    
		mem[    90] = 7'd29;    
		mem[    91] = 7'd30;    
		mem[    92] = 7'd29;    
		mem[    93] = 7'd30;    
		mem[    94] = 7'd29;    
		mem[    95] = 7'd30;    
		mem[    96] = 7'd29;    
		mem[    97] = 7'd29;    
		mem[    98] = 7'd30;    
		mem[    99] = 7'd29;    
		mem[   100] = 7'd30;    
		mem[   101] = 7'd29;    
		mem[   102] = 7'd30;    
		mem[   103] = 7'd29;    
		mem[   104] = 7'd29;    
		mem[   105] = 7'd30;    
		mem[   106] = 7'd29;    
		mem[   107] = 7'd30;    
		mem[   108] = 7'd29;    
		mem[   109] = 7'd30;    
		mem[   110] = 7'd29;    
		mem[   111] = 7'd30;    
		mem[   112] = 7'd29;    
		mem[   113] = 7'd29;    
		mem[   114] = 7'd30;    
		mem[   115] = 7'd29;    
		mem[   116] = 7'd30;    
		mem[   117] = 7'd29;    
		mem[   118] = 7'd30;    
		mem[   119] = 7'd29;    
		mem[   120] = 7'd30;    
		mem[   121] = 7'd29;    
		mem[   122] = 7'd29;    
		mem[   123] = 7'd30;    
		mem[   124] = 7'd29;    
		mem[   125] = 7'd59;    
		mem[   126] = 7'd29;    
		mem[   127] = 7'd30;    
		mem[   128] = 7'd29;    
		mem[   129] = 7'd30;    
		mem[   130] = 7'd30;    
		mem[   131] = 7'd29;    
		mem[   132] = 7'd29;    
		mem[   133] = 7'd30;    
		mem[   134] = 7'd29;    
		mem[   135] = 7'd30;    
		mem[   136] = 7'd6;    
		mem[   137] = 7'd8;    
		mem[   138] = 7'd45;    
		mem[   139] = 7'd29;    
		mem[   140] = 7'd29;    
		mem[   141] = 7'd30;    
		mem[   142] = 7'd29;    
		mem[   143] = 7'd29;    
		mem[   144] = 7'd30;    
		mem[   145] = 7'd29;    
		mem[   146] = 7'd29;    
		mem[   147] = 7'd30;    
		mem[   148] = 7'd29;    
		mem[   149] = 7'd30;    
		mem[   150] = 7'd29;    
		mem[   151] = 7'd30;    
		mem[   152] = 7'd29;    
		mem[   153] = 7'd30;    
		mem[   154] = 7'd29;    
		mem[   155] = 7'd30;    
		mem[   156] = 7'd29;    
		mem[   157] = 7'd29;    
		mem[   158] = 7'd30;    
		mem[   159] = 7'd29;    
		mem[   160] = 7'd30;    
		mem[   161] = 7'd29;    
		mem[   162] = 7'd30;    
		mem[   163] = 7'd29;    
		mem[   164] = 7'd29;    
		mem[   165] = 7'd30;    
		mem[   166] = 7'd29;    
		mem[   167] = 7'd30;    
		mem[   168] = 7'd29;    
		mem[   169] = 7'd30;    
		mem[   170] = 7'd29;    
		mem[   171] = 7'd30;    
		mem[   172] = 7'd29;    
		mem[   173] = 7'd30;    
		mem[   174] = 7'd29;    
		mem[   175] = 7'd30;    
		mem[   176] = 7'd29;    
		mem[   177] = 7'd29;    
		mem[   178] = 7'd30;    
		mem[   179] = 7'd29;    
		mem[   180] = 7'd30;    
		mem[   181] = 7'd29;    
		mem[   182] = 7'd29;    
		mem[   183] = 7'd30;    
		mem[   184] = 7'd29;    
		mem[   185] = 7'd30;    
		mem[   186] = 7'd29;    
		mem[   187] = 7'd30;    
		mem[   188] = 7'd29;    
		mem[   189] = 7'd30;    
		mem[   190] = 7'd29;    
		mem[   191] = 7'd30;    
		mem[   192] = 7'd29;    
		mem[   193] = 7'd29;    
		mem[   194] = 7'd30;    
		mem[   195] = 7'd29;    
		mem[   196] = 7'd30;    
		mem[   197] = 7'd29;    
		mem[   198] = 7'd29;    
		mem[   199] = 7'd30;    
		mem[   200] = 7'd29;    
		mem[   201] = 7'd30;    
		mem[   202] = 7'd29;    
		mem[   203] = 7'd30;    
		mem[   204] = 7'd29;    
		mem[   205] = 7'd30;    
		mem[   206] = 7'd29;    
		mem[   207] = 7'd30;    
		mem[   208] = 7'd29;    
		mem[   209] = 7'd29;    
		mem[   210] = 7'd30;    
		mem[   211] = 7'd29;    
		mem[   212] = 7'd30;    
		mem[   213] = 7'd29;    
		mem[   214] = 7'd29;    
		mem[   215] = 7'd30;    
		mem[   216] = 7'd29;    
		mem[   217] = 7'd30;    
		mem[   218] = 7'd29;    
		mem[   219] = 7'd30;    
		mem[   220] = 7'd29;    
		mem[   221] = 7'd30;    
		mem[   222] = 7'd29;    
		mem[   223] = 7'd30;    
		mem[   224] = 7'd29;    
		mem[   225] = 7'd30;    
		mem[   226] = 7'd29;    
		mem[   227] = 7'd29;    
		mem[   228] = 7'd30;    
		mem[   229] = 7'd29;    
		mem[   230] = 7'd30;    
		mem[   231] = 7'd29;    
		mem[   232] = 7'd29;    
		mem[   233] = 7'd30;    
		mem[   234] = 7'd29;    
		mem[   235] = 7'd30;    
		mem[   236] = 7'd29;    
		mem[   237] = 7'd30;    
		mem[   238] = 7'd29;    
		mem[   239] = 7'd30;    
		mem[   240] = 7'd29;    
		mem[   241] = 7'd29;    
		mem[   242] = 7'd30;    
		mem[   243] = 7'd29;    
		mem[   244] = 7'd30;    
		mem[   245] = 7'd29;    
		mem[   246] = 7'd30;    
		mem[   247] = 7'd29;    
		mem[   248] = 7'd29;    
		mem[   249] = 7'd30;    
		mem[   250] = 7'd29;    
		mem[   251] = 7'd30;    
		mem[   252] = 7'd29;    
		mem[   253] = 7'd30;    
		mem[   254] = 7'd29;    
		mem[   255] = 7'd30;    
		mem[   256] = 7'd29;    
		mem[   257] = 7'd30;    
		mem[   258] = 7'd29;    
		mem[   259] = 7'd29;    
		mem[   260] = 7'd29;    
		mem[   261] = 7'd60;    
		mem[   262] = 7'd29;    
		mem[   263] = 7'd30;    
		mem[   264] = 7'd29;    
		mem[   265] = 7'd29;    
		mem[   266] = 7'd30;    
		mem[   267] = 7'd29;    
		mem[   268] = 7'd30;    
		mem[   269] = 7'd29;    
		mem[   270] = 7'd30;    
		mem[   271] = 7'd29;    
		mem[   272] = 7'd59;    
		mem[   273] = 7'd59;    
		mem[   274] = 7'd59;    
		mem[   275] = 7'd59;    
		mem[   276] = 7'd29;    
		mem[   277] = 7'd30;    
		mem[   278] = 7'd61;    
		mem[   279] = 7'd29;    
		mem[   280] = 7'd44;    
		mem[   281] = 7'd13;    
		mem[   282] = 7'd17;    
		mem[   283] = 7'd28;    
		mem[   284] = 7'd29;    
		mem[   285] = 7'd29;    
		mem[   286] = 7'd30;    
		mem[   287] = 7'd29;    
		mem[   288] = 7'd30;    
		mem[   289] = 7'd29;    
		mem[   290] = 7'd29;    
		mem[   291] = 7'd30;    
		mem[   292] = 7'd29;    
		mem[   293] = 7'd30;    
		mem[   294] = 7'd29;    
		mem[   295] = 7'd29;    
		mem[   296] = 7'd30;    
		mem[   297] = 7'd29;    
		mem[   298] = 7'd30;    
		mem[   299] = 7'd29;    
		mem[   300] = 7'd30;    
		mem[   301] = 7'd29;    
		mem[   302] = 7'd30;    
		mem[   303] = 7'd29;    
		mem[   304] = 7'd29;    
		mem[   305] = 7'd30;    
		mem[   306] = 7'd29;    
		mem[   307] = 7'd30;    
		mem[   308] = 7'd29;    
		mem[   309] = 7'd30;    
		mem[   310] = 7'd29;    
		mem[   311] = 7'd30;    
		mem[   312] = 7'd29;    
		mem[   313] = 7'd30;    
		mem[   314] = 7'd29;    
		mem[   315] = 7'd29;    
		mem[   316] = 7'd30;    
		mem[   317] = 7'd29;    
		mem[   318] = 7'd30;    
		mem[   319] = 7'd29;    
		mem[   320] = 7'd30;    
		mem[   321] = 7'd29;    
		mem[   322] = 7'd30;    
		mem[   323] = 7'd29;    
		mem[   324] = 7'd30;    
		mem[   325] = 7'd29;    
		mem[   326] = 7'd29;    
		mem[   327] = 7'd30;    
		mem[   328] = 7'd29;    
		mem[   329] = 7'd30;    
		mem[   330] = 7'd29;    
		mem[   331] = 7'd30;    
		mem[   332] = 7'd29;    
		mem[   333] = 7'd29;    
		mem[   334] = 7'd30;    
		mem[   335] = 7'd29;    
		mem[   336] = 7'd30;    
		mem[   337] = 7'd29;    
		mem[   338] = 7'd30;    
		mem[   339] = 7'd29;    
		mem[   340] = 7'd30;    
		mem[   341] = 7'd29;    
		mem[   342] = 7'd29;    
		mem[   343] = 7'd30;    
		mem[   344] = 7'd29;    
		mem[   345] = 7'd30;    
		mem[   346] = 7'd29;    
		mem[   347] = 7'd30;    
		mem[   348] = 7'd29;    
		mem[   349] = 7'd30;    
		mem[   350] = 7'd29;    
		mem[   351] = 7'd29;    
		mem[   352] = 7'd30;    
		mem[   353] = 7'd29;    
		mem[   354] = 7'd30;    
		mem[   355] = 7'd29;    
		mem[   356] = 7'd30;    
		mem[   357] = 7'd29;    
		mem[   358] = 7'd30;    
		mem[   359] = 7'd29;    
		mem[   360] = 7'd30;    
		mem[   361] = 7'd29;    
		mem[   362] = 7'd29;    
		mem[   363] = 7'd30;    
		mem[   364] = 7'd29;    
		mem[   365] = 7'd30;    
		mem[   366] = 7'd29;    
		mem[   367] = 7'd29;    
		mem[   368] = 7'd30;    
		mem[   369] = 7'd29;    
		mem[   370] = 7'd30;    
		mem[   371] = 7'd29;    
		mem[   372] = 7'd30;    
		mem[   373] = 7'd29;    
		mem[   374] = 7'd30;    
		mem[   375] = 7'd29;    
		mem[   376] = 7'd29;    
		mem[   377] = 7'd30;    
		mem[   378] = 7'd29;    
		mem[   379] = 7'd30;    
		mem[   380] = 7'd29;    
		mem[   381] = 7'd30;    
		mem[   382] = 7'd29;    
		mem[   383] = 7'd29;    
		mem[   384] = 7'd30;    
		mem[   385] = 7'd29;    
		mem[   386] = 7'd30;    
		mem[   387] = 7'd29;    
		mem[   388] = 7'd30;    
		mem[   389] = 7'd29;    
		mem[   390] = 7'd30;    
		mem[   391] = 7'd29;    
		mem[   392] = 7'd29;    
		mem[   393] = 7'd30;    
		mem[   394] = 7'd29;    
		mem[   395] = 7'd30;    
		mem[   396] = 7'd29;    
		mem[   397] = 7'd30;    
		mem[   398] = 7'd29;    
		mem[   399] = 7'd30;    
		mem[   400] = 7'd29;    
		mem[   401] = 7'd29;    
		mem[   402] = 7'd30;    
		mem[   403] = 7'd29;    
		mem[   404] = 7'd59;    
		mem[   405] = 7'd29;    
		mem[   406] = 7'd30;    
		mem[   407] = 7'd29;    
		mem[   408] = 7'd30;    
		mem[   409] = 7'd30;    
		mem[   410] = 7'd29;    
		mem[   411] = 7'd29;    
		mem[   412] = 7'd30;    
		mem[   413] = 7'd29;    
		mem[   414] = 7'd30;    
		mem[   415] = 7'd6;    
		mem[   416] = 7'd8;    
		mem[   417] = 7'd45;    
		mem[   418] = 7'd29;    
		mem[   419] = 7'd29;    
		mem[   420] = 7'd30;    
		mem[   421] = 7'd29;    
		mem[   422] = 7'd29;    
		mem[   423] = 7'd30;    
		mem[   424] = 7'd29;    
		mem[   425] = 7'd29;    
		mem[   426] = 7'd30;    
		mem[   427] = 7'd29;    
		mem[   428] = 7'd30;    
		mem[   429] = 7'd29;    
		mem[   430] = 7'd30;    
		mem[   431] = 7'd29;    
		mem[   432] = 7'd30;    
		mem[   433] = 7'd29;    
		mem[   434] = 7'd30;    
		mem[   435] = 7'd29;    
		mem[   436] = 7'd29;    
		mem[   437] = 7'd30;    
		mem[   438] = 7'd29;    
		mem[   439] = 7'd30;    
		mem[   440] = 7'd29;    
		mem[   441] = 7'd30;    
		mem[   442] = 7'd29;    
		mem[   443] = 7'd29;    
		mem[   444] = 7'd30;    
		mem[   445] = 7'd29;    
		mem[   446] = 7'd30;    
		mem[   447] = 7'd29;    
		mem[   448] = 7'd30;    
		mem[   449] = 7'd29;    
		mem[   450] = 7'd30;    
		mem[   451] = 7'd29;    
		mem[   452] = 7'd30;    
		mem[   453] = 7'd29;    
		mem[   454] = 7'd30;    
		mem[   455] = 7'd29;    
		mem[   456] = 7'd29;    
		mem[   457] = 7'd30;    
		mem[   458] = 7'd29;    
		mem[   459] = 7'd30;    
		mem[   460] = 7'd29;    
		mem[   461] = 7'd29;    
		mem[   462] = 7'd30;    
		mem[   463] = 7'd29;    
		mem[   464] = 7'd30;    
		mem[   465] = 7'd29;    
		mem[   466] = 7'd30;    
		mem[   467] = 7'd29;    
		mem[   468] = 7'd30;    
		mem[   469] = 7'd29;    
		mem[   470] = 7'd30;    
		mem[   471] = 7'd29;    
		mem[   472] = 7'd29;    
		mem[   473] = 7'd30;    
		mem[   474] = 7'd29;    
		mem[   475] = 7'd30;    
		mem[   476] = 7'd29;    
		mem[   477] = 7'd29;    
		mem[   478] = 7'd30;    
		mem[   479] = 7'd29;    
		mem[   480] = 7'd30;    
		mem[   481] = 7'd29;    
		mem[   482] = 7'd30;    
		mem[   483] = 7'd29;    
		mem[   484] = 7'd30;    
		mem[   485] = 7'd29;    
		mem[   486] = 7'd30;    
		mem[   487] = 7'd29;    
		mem[   488] = 7'd29;    
		mem[   489] = 7'd30;    
		mem[   490] = 7'd29;    
		mem[   491] = 7'd30;    
		mem[   492] = 7'd29;    
		mem[   493] = 7'd29;    
		mem[   494] = 7'd30;    
		mem[   495] = 7'd29;    
		mem[   496] = 7'd30;    
		mem[   497] = 7'd29;    
		mem[   498] = 7'd30;    
		mem[   499] = 7'd29;    
		mem[   500] = 7'd30;    
		mem[   501] = 7'd29;    
		mem[   502] = 7'd30;    
		mem[   503] = 7'd29;    
		mem[   504] = 7'd30;    
		mem[   505] = 7'd29;    
		mem[   506] = 7'd29;    
		mem[   507] = 7'd30;    
		mem[   508] = 7'd29;    
		mem[   509] = 7'd30;    
		mem[   510] = 7'd29;    
		mem[   511] = 7'd29;    
		mem[   512] = 7'd30;    
		mem[   513] = 7'd29;    
		mem[   514] = 7'd30;    
		mem[   515] = 7'd29;    
		mem[   516] = 7'd30;    
		mem[   517] = 7'd29;    
		mem[   518] = 7'd30;    
		mem[   519] = 7'd29;    
		mem[   520] = 7'd29;    
		mem[   521] = 7'd30;    
		mem[   522] = 7'd29;    
		mem[   523] = 7'd30;    
		mem[   524] = 7'd29;    
		mem[   525] = 7'd30;    
		mem[   526] = 7'd29;    
		mem[   527] = 7'd29;    
		mem[   528] = 7'd30;    
		mem[   529] = 7'd29;    
		mem[   530] = 7'd30;    
		mem[   531] = 7'd29;    
		mem[   532] = 7'd30;    
		mem[   533] = 7'd29;    
		mem[   534] = 7'd30;    
		mem[   535] = 7'd29;    
		mem[   536] = 7'd30;    
		mem[   537] = 7'd29;    
		mem[   538] = 7'd29;    
		mem[   539] = 7'd29;    
		mem[   540] = 7'd60;    
		mem[   541] = 7'd29;    
		mem[   542] = 7'd30;    
		mem[   543] = 7'd29;    
		mem[   544] = 7'd29;    
		mem[   545] = 7'd30;    
		mem[   546] = 7'd29;    
		mem[   547] = 7'd30;    
		mem[   548] = 7'd29;    
		mem[   549] = 7'd30;    
		mem[   550] = 7'd29;    
		mem[   551] = 7'd59;    
		mem[   552] = 7'd59;    
		mem[   553] = 7'd59;    
		mem[   554] = 7'd59;    
		mem[   555] = 7'd29;    
		mem[   556] = 7'd30;    
		mem[   557] = 7'd61;    
		mem[   558] = 7'd29;    
		mem[   559] = 7'd44;    
		mem[   560] = 7'd13;    
		mem[   561] = 7'd17;    
		mem[   562] = 7'd28;    
		mem[   563] = 7'd29;    
		mem[   564] = 7'd29;    
		mem[   565] = 7'd30;    
		mem[   566] = 7'd29;    
		mem[   567] = 7'd30;    
		mem[   568] = 7'd29;    
		mem[   569] = 7'd29;    
		mem[   570] = 7'd30;    
		mem[   571] = 7'd29;    
		mem[   572] = 7'd30;    
		mem[   573] = 7'd29;    
		mem[   574] = 7'd29;    
		mem[   575] = 7'd30;    
		mem[   576] = 7'd29;    
		mem[   577] = 7'd30;    
		mem[   578] = 7'd29;    
		mem[   579] = 7'd30;    
		mem[   580] = 7'd29;    
		mem[   581] = 7'd30;    
		mem[   582] = 7'd29;    
		mem[   583] = 7'd29;    
		mem[   584] = 7'd30;    
		mem[   585] = 7'd29;    
		mem[   586] = 7'd30;    
		mem[   587] = 7'd29;    
		mem[   588] = 7'd30;    
		mem[   589] = 7'd29;    
		mem[   590] = 7'd30;    
		mem[   591] = 7'd29;    
		mem[   592] = 7'd30;    
		mem[   593] = 7'd29;    
		mem[   594] = 7'd29;    
		mem[   595] = 7'd30;    
		mem[   596] = 7'd29;    
		mem[   597] = 7'd30;    
		mem[   598] = 7'd29;    
		mem[   599] = 7'd30;    
		mem[   600] = 7'd29;    
		mem[   601] = 7'd30;    
		mem[   602] = 7'd29;    
		mem[   603] = 7'd30;    
		mem[   604] = 7'd29;    
		mem[   605] = 7'd29;    
		mem[   606] = 7'd30;    
		mem[   607] = 7'd29;    
		mem[   608] = 7'd30;    
		mem[   609] = 7'd29;    
		mem[   610] = 7'd30;    
		mem[   611] = 7'd29;    
		mem[   612] = 7'd29;    
		mem[   613] = 7'd30;    
		mem[   614] = 7'd29;    
		mem[   615] = 7'd30;    
		mem[   616] = 7'd29;    
		mem[   617] = 7'd30;    
		mem[   618] = 7'd29;    
		mem[   619] = 7'd30;    
		mem[   620] = 7'd29;    
		mem[   621] = 7'd29;    
		mem[   622] = 7'd30;    
		mem[   623] = 7'd29;    
		mem[   624] = 7'd30;    
		mem[   625] = 7'd29;    
		mem[   626] = 7'd30;    
		mem[   627] = 7'd29;    
		mem[   628] = 7'd30;    
		mem[   629] = 7'd29;    
		mem[   630] = 7'd29;    
		mem[   631] = 7'd30;    
		mem[   632] = 7'd29;    
		mem[   633] = 7'd30;    
		mem[   634] = 7'd29;    
		mem[   635] = 7'd30;    
		mem[   636] = 7'd29;    
		mem[   637] = 7'd30;    
		mem[   638] = 7'd29;    
		mem[   639] = 7'd30;    
		mem[   640] = 7'd29;    
		mem[   641] = 7'd29;    
		mem[   642] = 7'd30;    
		mem[   643] = 7'd29;    
		mem[   644] = 7'd30;    
		mem[   645] = 7'd29;    
		mem[   646] = 7'd29;    
		mem[   647] = 7'd30;    
		mem[   648] = 7'd29;    
		mem[   649] = 7'd30;    
		mem[   650] = 7'd29;    
		mem[   651] = 7'd30;    
		mem[   652] = 7'd29;    
		mem[   653] = 7'd30;    
		mem[   654] = 7'd29;    
		mem[   655] = 7'd29;    
		mem[   656] = 7'd30;    
		mem[   657] = 7'd29;    
		mem[   658] = 7'd30;    
		mem[   659] = 7'd29;    
		mem[   660] = 7'd30;    
		mem[   661] = 7'd29;    
		mem[   662] = 7'd29;    
		mem[   663] = 7'd30;    
		mem[   664] = 7'd29;    
		mem[   665] = 7'd30;    
		mem[   666] = 7'd29;    
		mem[   667] = 7'd30;    
		mem[   668] = 7'd29;    
		mem[   669] = 7'd30;    
		mem[   670] = 7'd29;    
		mem[   671] = 7'd29;    
		mem[   672] = 7'd30;    
		mem[   673] = 7'd29;    
		mem[   674] = 7'd30;    
		mem[   675] = 7'd29;    
		mem[   676] = 7'd30;    
		mem[   677] = 7'd29;    
		mem[   678] = 7'd30;    
		mem[   679] = 7'd29;    
		mem[   680] = 7'd29;    
		mem[   681] = 7'd30;    
		mem[   682] = 7'd29;    
		mem[   683] = 7'd59;    
		mem[   684] = 7'd29;    
		mem[   685] = 7'd30;    
		mem[   686] = 7'd29;    
		mem[   687] = 7'd30;    
		mem[   688] = 7'd30;    
		mem[   689] = 7'd29;    
		mem[   690] = 7'd29;    
		mem[   691] = 7'd30;    
		mem[   692] = 7'd29;    
		mem[   693] = 7'd30;    
		mem[   694] = 7'd6;    
		mem[   695] = 7'd8;    
		mem[   696] = 7'd45;    
		mem[   697] = 7'd29;    
		mem[   698] = 7'd29;    
		mem[   699] = 7'd30;    
		mem[   700] = 7'd29;    
		mem[   701] = 7'd29;    
		mem[   702] = 7'd30;    
		mem[   703] = 7'd29;    
		mem[   704] = 7'd29;    
		mem[   705] = 7'd30;    
		mem[   706] = 7'd29;    
		mem[   707] = 7'd30;    
		mem[   708] = 7'd29;    
		mem[   709] = 7'd30;    
		mem[   710] = 7'd29;    
		mem[   711] = 7'd30;    
		mem[   712] = 7'd29;    
		mem[   713] = 7'd30;    
		mem[   714] = 7'd29;    
		mem[   715] = 7'd29;    
		mem[   716] = 7'd30;    
		mem[   717] = 7'd29;    
		mem[   718] = 7'd30;    
		mem[   719] = 7'd29;    
		mem[   720] = 7'd30;    
		mem[   721] = 7'd29;    
		mem[   722] = 7'd29;    
		mem[   723] = 7'd30;    
		mem[   724] = 7'd29;    
		mem[   725] = 7'd30;    
		mem[   726] = 7'd29;    
		mem[   727] = 7'd30;    
		mem[   728] = 7'd29;    
		mem[   729] = 7'd30;    
		mem[   730] = 7'd29;    
		mem[   731] = 7'd30;    
		mem[   732] = 7'd29;    
		mem[   733] = 7'd30;    
		mem[   734] = 7'd29;    
		mem[   735] = 7'd29;    
		mem[   736] = 7'd30;    
		mem[   737] = 7'd29;    
		mem[   738] = 7'd30;    
		mem[   739] = 7'd29;    
		mem[   740] = 7'd29;    
		mem[   741] = 7'd30;    
		mem[   742] = 7'd29;    
		mem[   743] = 7'd30;    
		mem[   744] = 7'd29;    
		mem[   745] = 7'd30;    
		mem[   746] = 7'd29;    
		mem[   747] = 7'd30;    
		mem[   748] = 7'd29;    
		mem[   749] = 7'd30;    
		mem[   750] = 7'd29;    
		mem[   751] = 7'd29;    
		mem[   752] = 7'd30;    
		mem[   753] = 7'd29;    
		mem[   754] = 7'd30;    
		mem[   755] = 7'd29;    
		mem[   756] = 7'd29;    
		mem[   757] = 7'd30;    
		mem[   758] = 7'd29;    
		mem[   759] = 7'd30;    
		mem[   760] = 7'd29;    
		mem[   761] = 7'd30;    
		mem[   762] = 7'd29;    
		mem[   763] = 7'd30;    
		mem[   764] = 7'd29;    
		mem[   765] = 7'd30;    
		mem[   766] = 7'd29;    
		mem[   767] = 7'd29;    
		mem[   768] = 7'd30;    
		mem[   769] = 7'd29;    
		mem[   770] = 7'd30;    
		mem[   771] = 7'd29;    
		mem[   772] = 7'd29;    
		mem[   773] = 7'd30;    
		mem[   774] = 7'd29;    
		mem[   775] = 7'd30;    
		mem[   776] = 7'd29;    
		mem[   777] = 7'd30;    
		mem[   778] = 7'd29;    
		mem[   779] = 7'd30;    
		mem[   780] = 7'd29;    
		mem[   781] = 7'd30;    
		mem[   782] = 7'd29;    
		mem[   783] = 7'd30;    
		mem[   784] = 7'd29;    
		mem[   785] = 7'd29;    
		mem[   786] = 7'd30;    
		mem[   787] = 7'd29;    
		mem[   788] = 7'd30;    
		mem[   789] = 7'd29;    
		mem[   790] = 7'd29;    
		mem[   791] = 7'd30;    
		mem[   792] = 7'd29;    
		mem[   793] = 7'd30;    
		mem[   794] = 7'd29;    
		mem[   795] = 7'd30;    
		mem[   796] = 7'd29;    
		mem[   797] = 7'd30;    
		mem[   798] = 7'd29;    
		mem[   799] = 7'd29;    
		mem[   800] = 7'd30;    
		mem[   801] = 7'd29;    
		mem[   802] = 7'd30;    
		mem[   803] = 7'd29;    
		mem[   804] = 7'd30;    
		mem[   805] = 7'd29;    
		mem[   806] = 7'd29;    
		mem[   807] = 7'd30;    
		mem[   808] = 7'd29;    
		mem[   809] = 7'd30;    
		mem[   810] = 7'd29;    
		mem[   811] = 7'd30;    
		mem[   812] = 7'd29;    
		mem[   813] = 7'd30;    
		mem[   814] = 7'd29;    
		mem[   815] = 7'd30;    
		mem[   816] = 7'd29;    
		mem[   817] = 7'd29;    
		mem[   818] = 7'd29;    
		mem[   819] = 7'd60;    
		mem[   820] = 7'd29;    
		mem[   821] = 7'd30;    
		mem[   822] = 7'd29;    
		mem[   823] = 7'd29;    
		mem[   824] = 7'd30;    
		mem[   825] = 7'd29;    
		mem[   826] = 7'd30;    
		mem[   827] = 7'd29;    
		mem[   828] = 7'd30;    
		mem[   829] = 7'd29;    
		mem[   830] = 7'd59;    
		mem[   831] = 7'd59;    
		mem[   832] = 7'd59;    
		mem[   833] = 7'd59;    
		mem[   834] = 7'd29;    
		mem[   835] = 7'd30;    
		mem[   836] = 7'd61;    
		mem[   837] = 7'd29;    
		mem[   838] = 7'd44;    
		mem[   839] = 7'd13;    
		mem[   840] = 7'd17;    
		mem[   841] = 7'd28;    
		mem[   842] = 7'd29;    
		mem[   843] = 7'd29;    
		mem[   844] = 7'd30;    
		mem[   845] = 7'd29;    
		mem[   846] = 7'd30;    
		mem[   847] = 7'd29;    
		mem[   848] = 7'd29;    
		mem[   849] = 7'd30;    
		mem[   850] = 7'd29;    
		mem[   851] = 7'd30;    
		mem[   852] = 7'd29;    
		mem[   853] = 7'd29;    
		mem[   854] = 7'd30;    
		mem[   855] = 7'd29;    
		mem[   856] = 7'd30;    
		mem[   857] = 7'd29;    
		mem[   858] = 7'd30;    
		mem[   859] = 7'd29;    
		mem[   860] = 7'd30;    
		mem[   861] = 7'd29;    
		mem[   862] = 7'd29;    
		mem[   863] = 7'd30;    
		mem[   864] = 7'd29;    
		mem[   865] = 7'd30;    
		mem[   866] = 7'd29;    
		mem[   867] = 7'd30;    
		mem[   868] = 7'd29;    
		mem[   869] = 7'd30;    
		mem[   870] = 7'd29;    
		mem[   871] = 7'd30;    
		mem[   872] = 7'd29;    
		mem[   873] = 7'd29;    
		mem[   874] = 7'd30;    
		mem[   875] = 7'd29;    
		mem[   876] = 7'd30;    
		mem[   877] = 7'd29;    
		mem[   878] = 7'd30;    
		mem[   879] = 7'd29;    
		mem[   880] = 7'd30;    
		mem[   881] = 7'd29;    
		mem[   882] = 7'd30;    
		mem[   883] = 7'd29;    
		mem[   884] = 7'd29;    
		mem[   885] = 7'd30;    
		mem[   886] = 7'd29;    
		mem[   887] = 7'd30;    
		mem[   888] = 7'd29;    
		mem[   889] = 7'd30;    
		mem[   890] = 7'd29;    
		mem[   891] = 7'd29;    
		mem[   892] = 7'd30;    
		mem[   893] = 7'd29;    
		mem[   894] = 7'd30;    
		mem[   895] = 7'd29;    
		mem[   896] = 7'd30;    
		mem[   897] = 7'd29;    
		mem[   898] = 7'd30;    
		mem[   899] = 7'd29;    
		mem[   900] = 7'd29;    
		mem[   901] = 7'd30;    
		mem[   902] = 7'd29;    
		mem[   903] = 7'd30;    
		mem[   904] = 7'd29;    
		mem[   905] = 7'd30;    
		mem[   906] = 7'd29;    
		mem[   907] = 7'd30;    
		mem[   908] = 7'd29;    
		mem[   909] = 7'd29;    
		mem[   910] = 7'd30;    
		mem[   911] = 7'd29;    
		mem[   912] = 7'd30;    
		mem[   913] = 7'd29;    
		mem[   914] = 7'd30;    
		mem[   915] = 7'd29;    
		mem[   916] = 7'd30;    
		mem[   917] = 7'd29;    
		mem[   918] = 7'd30;    
		mem[   919] = 7'd29;    
		mem[   920] = 7'd29;    
		mem[   921] = 7'd30;    
		mem[   922] = 7'd29;    
		mem[   923] = 7'd30;    
		mem[   924] = 7'd29;    
		mem[   925] = 7'd29;    
		mem[   926] = 7'd30;    
		mem[   927] = 7'd29;    
		mem[   928] = 7'd30;    
		mem[   929] = 7'd29;    
		mem[   930] = 7'd30;    
		mem[   931] = 7'd29;    
		mem[   932] = 7'd30;    
		mem[   933] = 7'd29;    
		mem[   934] = 7'd29;    
		mem[   935] = 7'd30;    
		mem[   936] = 7'd29;    
		mem[   937] = 7'd30;    
		mem[   938] = 7'd29;    
		mem[   939] = 7'd30;    
		mem[   940] = 7'd29;    
		mem[   941] = 7'd29;    
		mem[   942] = 7'd30;    
		mem[   943] = 7'd29;    
		mem[   944] = 7'd30;    
		mem[   945] = 7'd29;    
		mem[   946] = 7'd30;    
		mem[   947] = 7'd29;    
		mem[   948] = 7'd30;    
		mem[   949] = 7'd29;    
		mem[   950] = 7'd29;    
		mem[   951] = 7'd30;    
		mem[   952] = 7'd29;    
		mem[   953] = 7'd30;    
		mem[   954] = 7'd29;    
		mem[   955] = 7'd30;    
		mem[   956] = 7'd29;    
		mem[   957] = 7'd30;    
		mem[   958] = 7'd29;    
		mem[   959] = 7'd29;    
		mem[   960] = 7'd30;    
		mem[   961] = 7'd29;    
		mem[   962] = 7'd59;    
		mem[   963] = 7'd29;    
		mem[   964] = 7'd30;    
		mem[   965] = 7'd29;    
		mem[   966] = 7'd30;    
		mem[   967] = 7'd30;    
		mem[   968] = 7'd29;    
		mem[   969] = 7'd29;    
		mem[   970] = 7'd30;    
		mem[   971] = 7'd29;    
		mem[   972] = 7'd30;    
		mem[   973] = 7'd6;    
		mem[   974] = 7'd8;    
		mem[   975] = 7'd45;    
		mem[   976] = 7'd29;    
		mem[   977] = 7'd29;    
		mem[   978] = 7'd30;    
		mem[   979] = 7'd29;    
		mem[   980] = 7'd29;    
		mem[   981] = 7'd30;    
		mem[   982] = 7'd29;    
		mem[   983] = 7'd29;    
		mem[   984] = 7'd30;    
		mem[   985] = 7'd29;    
		mem[   986] = 7'd30;    
		mem[   987] = 7'd29;    
		mem[   988] = 7'd30;    
		mem[   989] = 7'd29;    
		mem[   990] = 7'd30;    
		mem[   991] = 7'd29;    
		mem[   992] = 7'd30;    
		mem[   993] = 7'd29;    
		mem[   994] = 7'd29;    
		mem[   995] = 7'd30;    
		mem[   996] = 7'd29;    
		mem[   997] = 7'd30;    
		mem[   998] = 7'd29;    
		mem[   999] = 7'd30;    
		mem[  1000] = 7'd29;    
		mem[  1001] = 7'd29;    
		mem[  1002] = 7'd30;    
		mem[  1003] = 7'd29;    
		mem[  1004] = 7'd30;    
		mem[  1005] = 7'd29;    
		mem[  1006] = 7'd30;    
		mem[  1007] = 7'd29;    
		mem[  1008] = 7'd30;    
		mem[  1009] = 7'd29;    
		mem[  1010] = 7'd30;    
		mem[  1011] = 7'd29;    
		mem[  1012] = 7'd30;    
		mem[  1013] = 7'd29;    
		mem[  1014] = 7'd29;    
		mem[  1015] = 7'd30;    
		mem[  1016] = 7'd29;    
		mem[  1017] = 7'd30;    
		mem[  1018] = 7'd29;    
		mem[  1019] = 7'd29;    
		mem[  1020] = 7'd30;    
		mem[  1021] = 7'd29;    
		mem[  1022] = 7'd30;    
		mem[  1023] = 7'd29;    
		mem[  1024] = 7'd30;    
		mem[  1025] = 7'd29;    
		mem[  1026] = 7'd30;    
		mem[  1027] = 7'd29;    
		mem[  1028] = 7'd30;    
		mem[  1029] = 7'd29;    
		mem[  1030] = 7'd29;    
		mem[  1031] = 7'd30;    
		mem[  1032] = 7'd29;    
		mem[  1033] = 7'd30;    
		mem[  1034] = 7'd29;    
		mem[  1035] = 7'd29;    
		mem[  1036] = 7'd30;    
		mem[  1037] = 7'd29;    
		mem[  1038] = 7'd30;    
		mem[  1039] = 7'd29;    
		mem[  1040] = 7'd30;    
		mem[  1041] = 7'd29;    
		mem[  1042] = 7'd30;    
		mem[  1043] = 7'd29;    
		mem[  1044] = 7'd30;    
		mem[  1045] = 7'd29;    
		mem[  1046] = 7'd29;    
		mem[  1047] = 7'd30;    
		mem[  1048] = 7'd29;    
		mem[  1049] = 7'd30;    
		mem[  1050] = 7'd29;    
		mem[  1051] = 7'd29;    
		mem[  1052] = 7'd30;    
		mem[  1053] = 7'd29;    
		mem[  1054] = 7'd30;    
		mem[  1055] = 7'd29;    
		mem[  1056] = 7'd30;    
		mem[  1057] = 7'd29;    
		mem[  1058] = 7'd30;    
		mem[  1059] = 7'd29;    
		mem[  1060] = 7'd30;    
		mem[  1061] = 7'd29;    
		mem[  1062] = 7'd30;    
		mem[  1063] = 7'd29;    
		mem[  1064] = 7'd29;    
		mem[  1065] = 7'd30;    
		mem[  1066] = 7'd29;    
		mem[  1067] = 7'd30;    
		mem[  1068] = 7'd29;    
		mem[  1069] = 7'd29;    
		mem[  1070] = 7'd30;    
		mem[  1071] = 7'd29;    
		mem[  1072] = 7'd30;    
		mem[  1073] = 7'd29;    
		mem[  1074] = 7'd30;    
		mem[  1075] = 7'd29;    
		mem[  1076] = 7'd30;    
		mem[  1077] = 7'd29;    
		mem[  1078] = 7'd29;    
		mem[  1079] = 7'd30;    
		mem[  1080] = 7'd29;    
		mem[  1081] = 7'd30;    
		mem[  1082] = 7'd29;    
		mem[  1083] = 7'd30;    
		mem[  1084] = 7'd29;    
		mem[  1085] = 7'd29;    
		mem[  1086] = 7'd30;    
		mem[  1087] = 7'd29;    
		mem[  1088] = 7'd30;    
		mem[  1089] = 7'd29;    
		mem[  1090] = 7'd30;    
		mem[  1091] = 7'd29;    
		mem[  1092] = 7'd30;    
		mem[  1093] = 7'd29;    
		mem[  1094] = 7'd30;    
		mem[  1095] = 7'd29;    
		mem[  1096] = 7'd29;    
		mem[  1097] = 7'd29;    
		mem[  1098] = 7'd60;    
		mem[  1099] = 7'd29;    
		mem[  1100] = 7'd30;    
		mem[  1101] = 7'd29;    
		mem[  1102] = 7'd29;    
		mem[  1103] = 7'd30;    
		mem[  1104] = 7'd29;    
		mem[  1105] = 7'd30;    
		mem[  1106] = 7'd29;    
		mem[  1107] = 7'd30;    
		mem[  1108] = 7'd29;    
		mem[  1109] = 7'd59;    
		mem[  1110] = 7'd59;    
		mem[  1111] = 7'd59;    
		mem[  1112] = 7'd59;    
		mem[  1113] = 7'd29;    
		mem[  1114] = 7'd30;    
		mem[  1115] = 7'd61;    
		mem[  1116] = 7'd29;    
		mem[  1117] = 7'd44;    
		mem[  1118] = 7'd13;    
		mem[  1119] = 7'd17;    
		mem[  1120] = 7'd28;    
		mem[  1121] = 7'd29;    
		mem[  1122] = 7'd29;    
		mem[  1123] = 7'd30;    
		mem[  1124] = 7'd29;    
		mem[  1125] = 7'd30;    
		mem[  1126] = 7'd29;    
		mem[  1127] = 7'd29;    
		mem[  1128] = 7'd30;    
		mem[  1129] = 7'd29;    
		mem[  1130] = 7'd30;    
		mem[  1131] = 7'd29;    
		mem[  1132] = 7'd29;    
		mem[  1133] = 7'd30;    
		mem[  1134] = 7'd29;    
		mem[  1135] = 7'd30;    
		mem[  1136] = 7'd29;    
		mem[  1137] = 7'd30;    
		mem[  1138] = 7'd29;    
		mem[  1139] = 7'd30;    
		mem[  1140] = 7'd29;    
		mem[  1141] = 7'd29;    
		mem[  1142] = 7'd30;    
		mem[  1143] = 7'd29;    
		mem[  1144] = 7'd30;    
		mem[  1145] = 7'd29;    
		mem[  1146] = 7'd30;    
		mem[  1147] = 7'd29;    
		mem[  1148] = 7'd30;    
		mem[  1149] = 7'd29;    
		mem[  1150] = 7'd30;    
		mem[  1151] = 7'd29;    
		mem[  1152] = 7'd29;    
		mem[  1153] = 7'd30;    
		mem[  1154] = 7'd29;    
		mem[  1155] = 7'd30;    
		mem[  1156] = 7'd29;    
		mem[  1157] = 7'd30;    
		mem[  1158] = 7'd29;    
		mem[  1159] = 7'd30;    
		mem[  1160] = 7'd29;    
		mem[  1161] = 7'd30;    
		mem[  1162] = 7'd29;    
		mem[  1163] = 7'd29;    
		mem[  1164] = 7'd30;    
		mem[  1165] = 7'd29;    
		mem[  1166] = 7'd30;    
		mem[  1167] = 7'd29;    
		mem[  1168] = 7'd30;    
		mem[  1169] = 7'd29;    
		mem[  1170] = 7'd29;    
		mem[  1171] = 7'd30;    
		mem[  1172] = 7'd29;    
		mem[  1173] = 7'd30;    
		mem[  1174] = 7'd29;    
		mem[  1175] = 7'd30;    
		mem[  1176] = 7'd29;    
		mem[  1177] = 7'd30;    
		mem[  1178] = 7'd29;    
		mem[  1179] = 7'd29;    
		mem[  1180] = 7'd30;    
		mem[  1181] = 7'd29;    
		mem[  1182] = 7'd30;    
		mem[  1183] = 7'd29;    
		mem[  1184] = 7'd30;    
		mem[  1185] = 7'd29;    
		mem[  1186] = 7'd30;    
		mem[  1187] = 7'd29;    
		mem[  1188] = 7'd29;    
		mem[  1189] = 7'd30;    
		mem[  1190] = 7'd29;    
		mem[  1191] = 7'd30;    
		mem[  1192] = 7'd29;    
		mem[  1193] = 7'd30;    
		mem[  1194] = 7'd29;    
		mem[  1195] = 7'd30;    
		mem[  1196] = 7'd29;    
		mem[  1197] = 7'd30;    
		mem[  1198] = 7'd29;    
		mem[  1199] = 7'd29;    
		mem[  1200] = 7'd30;    
		mem[  1201] = 7'd29;    
		mem[  1202] = 7'd30;    
		mem[  1203] = 7'd29;    
		mem[  1204] = 7'd29;    
		mem[  1205] = 7'd30;    
		mem[  1206] = 7'd29;    
		mem[  1207] = 7'd30;    
		mem[  1208] = 7'd29;    
		mem[  1209] = 7'd30;    
		mem[  1210] = 7'd29;    
		mem[  1211] = 7'd30;    
		mem[  1212] = 7'd29;    
		mem[  1213] = 7'd29;    
		mem[  1214] = 7'd30;    
		mem[  1215] = 7'd29;    
		mem[  1216] = 7'd30;    
		mem[  1217] = 7'd29;    
		mem[  1218] = 7'd30;    
		mem[  1219] = 7'd29;    
		mem[  1220] = 7'd29;    
		mem[  1221] = 7'd30;    
		mem[  1222] = 7'd29;    
		mem[  1223] = 7'd30;    
		mem[  1224] = 7'd29;    
		mem[  1225] = 7'd30;    
		mem[  1226] = 7'd29;    
		mem[  1227] = 7'd30;    
		mem[  1228] = 7'd29;    
		mem[  1229] = 7'd29;    
		mem[  1230] = 7'd30;    
		mem[  1231] = 7'd29;    
		mem[  1232] = 7'd30;    
		mem[  1233] = 7'd29;    
		mem[  1234] = 7'd30;    
		mem[  1235] = 7'd29;    
		mem[  1236] = 7'd30;    
		mem[  1237] = 7'd29;    
		mem[  1238] = 7'd29;    
		mem[  1239] = 7'd30;    
		mem[  1240] = 7'd29;    
		mem[  1241] = 7'd59;    
		mem[  1242] = 7'd29;    
		mem[  1243] = 7'd30;    
		mem[  1244] = 7'd29;    
		mem[  1245] = 7'd30;    
		mem[  1246] = 7'd30;    
		mem[  1247] = 7'd29;    
		mem[  1248] = 7'd29;    
		mem[  1249] = 7'd30;    
		mem[  1250] = 7'd29;    
		mem[  1251] = 7'd30;    
		mem[  1252] = 7'd6;    
		mem[  1253] = 7'd8;    
		mem[  1254] = 7'd45;    
		mem[  1255] = 7'd29;    
		mem[  1256] = 7'd29;    
		mem[  1257] = 7'd30;    
		mem[  1258] = 7'd29;    
		mem[  1259] = 7'd29;    
		mem[  1260] = 7'd30;    
		mem[  1261] = 7'd29;    
		mem[  1262] = 7'd29;    
		mem[  1263] = 7'd30;    
		mem[  1264] = 7'd29;    
		mem[  1265] = 7'd30;    
		mem[  1266] = 7'd29;    
		mem[  1267] = 7'd30;    
		mem[  1268] = 7'd29;    
		mem[  1269] = 7'd30;    
		mem[  1270] = 7'd29;    
		mem[  1271] = 7'd30;    
		mem[  1272] = 7'd29;    
		mem[  1273] = 7'd29;    
		mem[  1274] = 7'd30;    
		mem[  1275] = 7'd29;    
		mem[  1276] = 7'd30;    
		mem[  1277] = 7'd29;    
		mem[  1278] = 7'd30;    
		mem[  1279] = 7'd29;    
		mem[  1280] = 7'd29;    
		mem[  1281] = 7'd30;    
		mem[  1282] = 7'd29;    
		mem[  1283] = 7'd30;    
		mem[  1284] = 7'd29;    
		mem[  1285] = 7'd30;    
		mem[  1286] = 7'd29;    
		mem[  1287] = 7'd30;    
		mem[  1288] = 7'd29;    
		mem[  1289] = 7'd30;    
		mem[  1290] = 7'd29;    
		mem[  1291] = 7'd30;    
		mem[  1292] = 7'd29;    
		mem[  1293] = 7'd29;    
		mem[  1294] = 7'd30;    
		mem[  1295] = 7'd29;    
		mem[  1296] = 7'd30;    
		mem[  1297] = 7'd29;    
		mem[  1298] = 7'd29;    
		mem[  1299] = 7'd30;    
		mem[  1300] = 7'd29;    
		mem[  1301] = 7'd30;    
		mem[  1302] = 7'd29;    
		mem[  1303] = 7'd30;    
		mem[  1304] = 7'd29;    
		mem[  1305] = 7'd30;    
		mem[  1306] = 7'd29;    
		mem[  1307] = 7'd30;    
		mem[  1308] = 7'd29;    
		mem[  1309] = 7'd29;    
		mem[  1310] = 7'd30;    
		mem[  1311] = 7'd29;    
		mem[  1312] = 7'd30;    
		mem[  1313] = 7'd29;    
		mem[  1314] = 7'd29;    
		mem[  1315] = 7'd30;    
		mem[  1316] = 7'd29;    
		mem[  1317] = 7'd30;    
		mem[  1318] = 7'd29;    
		mem[  1319] = 7'd30;    
		mem[  1320] = 7'd29;    
		mem[  1321] = 7'd30;    
		mem[  1322] = 7'd29;    
		mem[  1323] = 7'd30;    
		mem[  1324] = 7'd29;    
		mem[  1325] = 7'd29;    
		mem[  1326] = 7'd30;    
		mem[  1327] = 7'd29;    
		mem[  1328] = 7'd30;    
		mem[  1329] = 7'd29;    
		mem[  1330] = 7'd29;    
		mem[  1331] = 7'd30;    
		mem[  1332] = 7'd29;    
		mem[  1333] = 7'd30;    
		mem[  1334] = 7'd29;    
		mem[  1335] = 7'd30;    
		mem[  1336] = 7'd29;    
		mem[  1337] = 7'd30;    
		mem[  1338] = 7'd29;    
		mem[  1339] = 7'd30;    
		mem[  1340] = 7'd29;    
		mem[  1341] = 7'd30;    
		mem[  1342] = 7'd29;    
		mem[  1343] = 7'd29;    
		mem[  1344] = 7'd30;    
		mem[  1345] = 7'd29;    
		mem[  1346] = 7'd30;    
		mem[  1347] = 7'd29;    
		mem[  1348] = 7'd29;    
		mem[  1349] = 7'd30;    
		mem[  1350] = 7'd29;    
		mem[  1351] = 7'd30;    
		mem[  1352] = 7'd29;    
		mem[  1353] = 7'd30;    
		mem[  1354] = 7'd29;    
		mem[  1355] = 7'd30;    
		mem[  1356] = 7'd29;    
		mem[  1357] = 7'd29;    
		mem[  1358] = 7'd30;    
		mem[  1359] = 7'd29;    
		mem[  1360] = 7'd30;    
		mem[  1361] = 7'd29;    
		mem[  1362] = 7'd30;    
		mem[  1363] = 7'd29;    
		mem[  1364] = 7'd29;    
		mem[  1365] = 7'd30;    
		mem[  1366] = 7'd29;    
		mem[  1367] = 7'd30;    
		mem[  1368] = 7'd29;    
		mem[  1369] = 7'd30;    
		mem[  1370] = 7'd29;    
		mem[  1371] = 7'd30;    
		mem[  1372] = 7'd29;    
		mem[  1373] = 7'd30;    
		mem[  1374] = 7'd29;    
		mem[  1375] = 7'd29;    
		mem[  1376] = 7'd29;    
		mem[  1377] = 7'd60;    
		mem[  1378] = 7'd29;    
		mem[  1379] = 7'd30;    
		mem[  1380] = 7'd29;    
		mem[  1381] = 7'd29;    
		mem[  1382] = 7'd30;    
		mem[  1383] = 7'd29;    
		mem[  1384] = 7'd30;    
		mem[  1385] = 7'd29;    
		mem[  1386] = 7'd30;    
		mem[  1387] = 7'd29;    
		mem[  1388] = 7'd59;    
		mem[  1389] = 7'd59;    
		mem[  1390] = 7'd59;    
		mem[  1391] = 7'd59;    
		mem[  1392] = 7'd29;    
		mem[  1393] = 7'd30;    
		mem[  1394] = 7'd59;     
	end
	
endmodule

