module pacman_intermission_converted2(in, out, clk); //ok
	 input [11:0] in;
	 input clk;
	 output reg [10:0] out;
	 
	 reg  [10:0] mem [0:2182];
	 always @(posedge clk) out  =  mem[ in ];
	 
	 initial begin
		mem[     0] = 11'd190;    
		mem[     1] = 11'd43;    
		mem[     2] = 11'd39;    
		mem[     3] = 11'd49;    
		mem[     4] = 11'd40;    
		mem[     5] = 11'd32;    
		mem[     6] = 11'd43;    
		mem[     7] = 11'd48;    
		mem[     8] = 11'd31;    
		mem[     9] = 11'd43;    
		mem[    10] = 11'd89;    
		mem[    11] = 11'd41;    
		mem[    12] = 11'd33;    
		mem[    13] = 11'd43;    
		mem[    14] = 11'd48;    
		mem[    15] = 11'd31;    
		mem[    16] = 11'd43;    
		mem[    17] = 11'd40;    
		mem[    18] = 11'd49;    
		mem[    19] = 11'd41;    
		mem[    20] = 11'd33;    
		mem[    21] = 11'd44;    
		mem[    22] = 11'd47;    
		mem[    23] = 11'd31;    
		mem[    24] = 11'd44;    
		mem[    25] = 11'd40;    
		mem[    26] = 11'd48;    
		mem[    27] = 11'd41;    
		mem[    28] = 11'd34;    
		mem[    29] = 11'd43;    
		mem[    30] = 11'd46;    
		mem[    31] = 11'd32;    
		mem[    32] = 11'd44;    
		mem[    33] = 11'd159;    
		mem[    34] = 11'd113;    
		mem[    35] = 11'd42;    
		mem[    36] = 11'd156;    
		mem[    37] = 11'd130;    
		mem[    38] = 11'd42;    
		mem[    39] = 11'd162;    
		mem[    40] = 11'd124;    
		mem[    41] = 11'd42;    
		mem[    42] = 11'd162;    
		mem[    43] = 11'd124;    
		mem[    44] = 11'd42;    
		mem[    45] = 11'd162;    
		mem[    46] = 11'd76;    
		mem[    47] = 11'd22;    
		mem[    48] = 11'd20;    
		mem[    49] = 11'd18;    
		mem[    50] = 11'd24;    
		mem[    51] = 11'd19;    
		mem[    52] = 11'd20;    
		mem[    53] = 11'd21;    
		mem[    54] = 11'd21;    
		mem[    55] = 11'd22;    
		mem[    56] = 11'd21;    
		mem[    57] = 11'd20;    
		mem[    58] = 11'd20;    
		mem[    59] = 11'd19;    
		mem[    60] = 11'd20;    
		mem[    61] = 11'd22;    
		mem[    62] = 11'd22;    
		mem[    63] = 11'd20;    
		mem[    64] = 11'd20;    
		mem[    65] = 11'd19;    
		mem[    66] = 11'd23;    
		mem[    67] = 11'd19;    
		mem[    68] = 11'd20;    
		mem[    69] = 11'd20;    
		mem[    70] = 11'd21;    
		mem[    71] = 11'd22;    
		mem[    72] = 11'd20;    
		mem[    73] = 11'd21;    
		mem[    74] = 11'd19;    
		mem[    75] = 11'd20;    
		mem[    76] = 11'd20;    
		mem[    77] = 11'd21;    
		mem[    78] = 11'd22;    
		mem[    79] = 11'd21;    
		mem[    80] = 11'd19;    
		mem[    81] = 11'd19;    
		mem[    82] = 11'd23;    
		mem[    83] = 11'd19;    
		mem[    84] = 11'd20;    
		mem[    85] = 11'd21;    
		mem[    86] = 11'd21;    
		mem[    87] = 11'd21;    
		mem[    88] = 11'd21;    
		mem[    89] = 11'd20;    
		mem[    90] = 11'd20;    
		mem[    91] = 11'd20;    
		mem[    92] = 11'd20;    
		mem[    93] = 11'd21;    
		mem[    94] = 11'd21;    
		mem[    95] = 11'd21;    
		mem[    96] = 11'd20;    
		mem[    97] = 11'd19;    
		mem[    98] = 11'd22;    
		mem[    99] = 11'd20;    
		mem[   100] = 11'd20;    
		mem[   101] = 11'd21;    
		mem[   102] = 11'd20;    
		mem[   103] = 11'd21;    
		mem[   104] = 11'd21;    
		mem[   105] = 11'd20;    
		mem[   106] = 11'd21;    
		mem[   107] = 11'd19;    
		mem[   108] = 11'd21;    
		mem[   109] = 11'd21;    
		mem[   110] = 11'd21;    
		mem[   111] = 11'd20;    
		mem[   112] = 11'd21;    
		mem[   113] = 11'd19;    
		mem[   114] = 11'd22;    
		mem[   115] = 11'd177;    
		mem[   116] = 11'd108;    
		mem[   117] = 11'd47;    
		mem[   118] = 11'd1146;    
		mem[   119] = 11'd27;    
		mem[   120] = 11'd27;    
		mem[   121] = 11'd27;    
		mem[   122] = 11'd27;    
		mem[   123] = 11'd28;    
		mem[   124] = 11'd27;    
		mem[   125] = 11'd27;    
		mem[   126] = 11'd27;    
		mem[   127] = 11'd28;    
		mem[   128] = 11'd27;    
		mem[   129] = 11'd27;    
		mem[   130] = 11'd28;    
		mem[   131] = 11'd27;    
		mem[   132] = 11'd27;    
		mem[   133] = 11'd27;    
		mem[   134] = 11'd28;    
		mem[   135] = 11'd27;    
		mem[   136] = 11'd27;    
		mem[   137] = 11'd28;    
		mem[   138] = 11'd27;    
		mem[   139] = 11'd27;    
		mem[   140] = 11'd27;    
		mem[   141] = 11'd28;    
		mem[   142] = 11'd27;    
		mem[   143] = 11'd28;    
		mem[   144] = 11'd27;    
		mem[   145] = 11'd27;    
		mem[   146] = 11'd27;    
		mem[   147] = 11'd28;    
		mem[   148] = 11'd27;    
		mem[   149] = 11'd27;    
		mem[   150] = 11'd28;    
		mem[   151] = 11'd27;    
		mem[   152] = 11'd27;    
		mem[   153] = 11'd28;    
		mem[   154] = 11'd27;    
		mem[   155] = 11'd27;    
		mem[   156] = 11'd28;    
		mem[   157] = 11'd27;    
		mem[   158] = 11'd27;    
		mem[   159] = 11'd27;    
		mem[   160] = 11'd28;    
		mem[   161] = 11'd27;    
		mem[   162] = 11'd27;    
		mem[   163] = 11'd28;    
		mem[   164] = 11'd27;    
		mem[   165] = 11'd27;    
		mem[   166] = 11'd28;    
		mem[   167] = 11'd27;    
		mem[   168] = 11'd27;    
		mem[   169] = 11'd27;    
		mem[   170] = 11'd28;    
		mem[   171] = 11'd27;    
		mem[   172] = 11'd1101;    
		mem[   173] = 11'd387;    
		mem[   174] = 11'd66;    
		mem[   175] = 11'd31;    
		mem[   176] = 11'd30;    
		mem[   177] = 11'd41;    
		mem[   178] = 11'd28;    
		mem[   179] = 11'd68;    
		mem[   180] = 11'd23;    
		mem[   181] = 11'd20;    
		mem[   182] = 11'd14;    
		mem[   183] = 11'd34;    
		mem[   184] = 11'd39;    
		mem[   185] = 11'd27;    
		mem[   186] = 11'd31;    
		mem[   187] = 11'd38;    
		mem[   188] = 11'd33;    
		mem[   189] = 11'd24;    
		mem[   190] = 11'd38;    
		mem[   191] = 11'd35;    
		mem[   192] = 11'd26;    
		mem[   193] = 11'd39;    
		mem[   194] = 11'd31;    
		mem[   195] = 11'd31;    
		mem[   196] = 11'd27;    
		mem[   197] = 11'd41;    
		mem[   198] = 11'd31;    
		mem[   199] = 11'd26;    
		mem[   200] = 11'd41;    
		mem[   201] = 11'd28;    
		mem[   202] = 11'd31;    
		mem[   203] = 11'd32;    
		mem[   204] = 11'd40;    
		mem[   205] = 11'd28;    
		mem[   206] = 11'd29;    
		mem[   207] = 11'd39;    
		mem[   208] = 11'd24;    
		mem[   209] = 11'd35;    
		mem[   210] = 11'd35;    
		mem[   211] = 11'd36;    
		mem[   212] = 11'd27;    
		mem[   213] = 11'd34;    
		mem[   214] = 11'd35;    
		mem[   215] = 11'd33;    
		mem[   216] = 11'd27;    
		mem[   217] = 11'd70;    
		mem[   218] = 11'd95;    
		mem[   219] = 11'd28;    
		mem[   220] = 11'd110;    
		mem[   221] = 11'd85;    
		mem[   222] = 11'd28;    
		mem[   223] = 11'd109;    
		mem[   224] = 11'd81;    
		mem[   225] = 11'd28;    
		mem[   226] = 11'd105;    
		mem[   227] = 11'd82;    
		mem[   228] = 11'd28;    
		mem[   229] = 11'd109;    
		mem[   230] = 11'd81;    
		mem[   231] = 11'd28;    
		mem[   232] = 11'd108;    
		mem[   233] = 11'd83;    
		mem[   234] = 11'd30;    
		mem[   235] = 11'd106;    
		mem[   236] = 11'd93;    
		mem[   237] = 11'd20;    
		mem[   238] = 11'd19;    
		mem[   239] = 11'd18;    
		mem[   240] = 11'd19;    
		mem[   241] = 11'd22;    
		mem[   242] = 11'd23;    
		mem[   243] = 11'd23;    
		mem[   244] = 11'd20;    
		mem[   245] = 11'd18;    
		mem[   246] = 11'd18;    
		mem[   247] = 11'd18;    
		mem[   248] = 11'd44;    
		mem[   249] = 11'd23;    
		mem[   250] = 11'd20;    
		mem[   251] = 11'd18;    
		mem[   252] = 11'd20;    
		mem[   253] = 11'd21;    
		mem[   254] = 11'd18;    
		mem[   255] = 11'd42;    
		mem[   256] = 11'd23;    
		mem[   257] = 11'd22;    
		mem[   258] = 11'd21;    
		mem[   259] = 11'd19;    
		mem[   260] = 11'd19;    
		mem[   261] = 11'd17;    
		mem[   262] = 11'd45;    
		mem[   263] = 11'd23;    
		mem[   264] = 11'd20;    
		mem[   265] = 11'd17;    
		mem[   266] = 11'd21;    
		mem[   267] = 11'd20;    
		mem[   268] = 11'd19;    
		mem[   269] = 11'd20;    
		mem[   270] = 11'd22;    
		mem[   271] = 11'd22;    
		mem[   272] = 11'd23;    
		mem[   273] = 11'd21;    
		mem[   274] = 11'd18;    
		mem[   275] = 11'd19;    
		mem[   276] = 11'd18;    
		mem[   277] = 11'd21;    
		mem[   278] = 11'd24;    
		mem[   279] = 11'd22;    
		mem[   280] = 11'd20;    
		mem[   281] = 11'd18;    
		mem[   282] = 11'd21;    
		mem[   283] = 11'd20;    
		mem[   284] = 11'd19;    
		mem[   285] = 11'd19;    
		mem[   286] = 11'd23;    
		mem[   287] = 11'd22;    
		mem[   288] = 11'd22;    
		mem[   289] = 11'd21;    
		mem[   290] = 11'd19;    
		mem[   291] = 11'd19;    
		mem[   292] = 11'd18;    
		mem[   293] = 11'd21;    
		mem[   294] = 11'd23;    
		mem[   295] = 11'd23;    
		mem[   296] = 11'd20;    
		mem[   297] = 11'd18;    
		mem[   298] = 11'd20;    
		mem[   299] = 11'd21;    
		mem[   300] = 11'd19;    
		mem[   301] = 11'd20;    
		mem[   302] = 11'd21;    
		mem[   303] = 11'd23;    
		mem[   304] = 11'd27;    
		mem[   305] = 11'd27;    
		mem[   306] = 11'd24;    
		mem[   307] = 11'd25;    
		mem[   308] = 11'd29;    
		mem[   309] = 11'd32;    
		mem[   310] = 11'd26;    
		mem[   311] = 11'd22;    
		mem[   312] = 11'd31;    
		mem[   313] = 11'd25;    
		mem[   314] = 11'd27;    
		mem[   315] = 11'd30;    
		mem[   316] = 11'd30;    
		mem[   317] = 11'd26;    
		mem[   318] = 11'd25;    
		mem[   319] = 11'd25;    
		mem[   320] = 11'd29;    
		mem[   321] = 11'd31;    
		mem[   322] = 11'd26;    
		mem[   323] = 11'd23;    
		mem[   324] = 11'd30;    
		mem[   325] = 11'd25;    
		mem[   326] = 11'd28;    
		mem[   327] = 11'd30;    
		mem[   328] = 11'd29;    
		mem[   329] = 11'd27;    
		mem[   330] = 11'd25;    
		mem[   331] = 11'd25;    
		mem[   332] = 11'd29;    
		mem[   333] = 11'd30;    
		mem[   334] = 11'd27;    
		mem[   335] = 11'd23;    
		mem[   336] = 11'd30;    
		mem[   337] = 11'd25;    
		mem[   338] = 11'd28;    
		mem[   339] = 11'd30;    
		mem[   340] = 11'd29;    
		mem[   341] = 11'd26;    
		mem[   342] = 11'd25;    
		mem[   343] = 11'd25;    
		mem[   344] = 11'd30;    
		mem[   345] = 11'd29;    
		mem[   346] = 11'd27;    
		mem[   347] = 11'd24;    
		mem[   348] = 11'd30;    
		mem[   349] = 11'd25;    
		mem[   350] = 11'd28;    
		mem[   351] = 11'd29;    
		mem[   352] = 11'd29;    
		mem[   353] = 11'd27;    
		mem[   354] = 11'd25;    
		mem[   355] = 11'd26;    
		mem[   356] = 11'd28;    
		mem[   357] = 11'd81;    
		mem[   358] = 11'd48;    
		mem[   359] = 11'd140;    
		mem[   360] = 11'd118;    
		mem[   361] = 11'd50;    
		mem[   362] = 11'd154;    
		mem[   363] = 11'd132;    
		mem[   364] = 11'd42;    
		mem[   365] = 11'd162;    
		mem[   366] = 11'd124;    
		mem[   367] = 11'd42;    
		mem[   368] = 11'd162;    
		mem[   369] = 11'd124;    
		mem[   370] = 11'd42;    
		mem[   371] = 11'd163;    
		mem[   372] = 11'd123;    
		mem[   373] = 11'd42;    
		mem[   374] = 11'd168;    
		mem[   375] = 11'd118;    
		mem[   376] = 11'd44;    
		mem[   377] = 11'd926;    
		mem[   378] = 11'd34;    
		mem[   379] = 11'd34;    
		mem[   380] = 11'd33;    
		mem[   381] = 11'd33;    
		mem[   382] = 11'd33;    
		mem[   383] = 11'd33;    
		mem[   384] = 11'd32;    
		mem[   385] = 11'd33;    
		mem[   386] = 11'd32;    
		mem[   387] = 11'd33;    
		mem[   388] = 11'd32;    
		mem[   389] = 11'd33;    
		mem[   390] = 11'd32;    
		mem[   391] = 11'd33;    
		mem[   392] = 11'd32;    
		mem[   393] = 11'd32;    
		mem[   394] = 11'd33;    
		mem[   395] = 11'd32;    
		mem[   396] = 11'd33;    
		mem[   397] = 11'd32;    
		mem[   398] = 11'd33;    
		mem[   399] = 11'd32;    
		mem[   400] = 11'd32;    
		mem[   401] = 11'd33;    
		mem[   402] = 11'd32;    
		mem[   403] = 11'd33;    
		mem[   404] = 11'd32;    
		mem[   405] = 11'd33;    
		mem[   406] = 11'd32;    
		mem[   407] = 11'd33;    
		mem[   408] = 11'd32;    
		mem[   409] = 11'd33;    
		mem[   410] = 11'd32;    
		mem[   411] = 11'd33;    
		mem[   412] = 11'd32;    
		mem[   413] = 11'd32;    
		mem[   414] = 11'd33;    
		mem[   415] = 11'd32;    
		mem[   416] = 11'd33;    
		mem[   417] = 11'd32;    
		mem[   418] = 11'd33;    
		mem[   419] = 11'd32;    
		mem[   420] = 11'd33;    
		mem[   421] = 11'd32;    
		mem[   422] = 11'd33;    
		mem[   423] = 11'd32;    
		mem[   424] = 11'd33;    
		mem[   425] = 11'd32;    
		mem[   426] = 11'd33;    
		mem[   427] = 11'd32;    
		mem[   428] = 11'd33;    
		mem[   429] = 11'd32;    
		mem[   430] = 11'd32;    
		mem[   431] = 11'd33;    
		mem[   432] = 11'd33;    
		mem[   433] = 11'd32;    
		mem[   434] = 11'd33;    
		mem[   435] = 11'd32;    
		mem[   436] = 11'd32;    
		mem[   437] = 11'd33;    
		mem[   438] = 11'd32;    
		mem[   439] = 11'd33;    
		mem[   440] = 11'd32;    
		mem[   441] = 11'd33;    
		mem[   442] = 11'd32;    
		mem[   443] = 11'd33;    
		mem[   444] = 11'd32;    
		mem[   445] = 11'd33;    
		mem[   446] = 11'd32;    
		mem[   447] = 11'd33;    
		mem[   448] = 11'd32;    
		mem[   449] = 11'd33;    
		mem[   450] = 11'd32;    
		mem[   451] = 11'd33;    
		mem[   452] = 11'd32;    
		mem[   453] = 11'd33;    
		mem[   454] = 11'd32;    
		mem[   455] = 11'd33;    
		mem[   456] = 11'd32;    
		mem[   457] = 11'd33;    
		mem[   458] = 11'd32;    
		mem[   459] = 11'd33;    
		mem[   460] = 11'd32;    
		mem[   461] = 11'd33;    
		mem[   462] = 11'd32;    
		mem[   463] = 11'd33;    
		mem[   464] = 11'd32;    
		mem[   465] = 11'd70;    
		mem[   466] = 11'd28;    
		mem[   467] = 11'd107;    
		mem[   468] = 11'd83;    
		mem[   469] = 11'd27;    
		mem[   470] = 11'd108;    
		mem[   471] = 11'd83;    
		mem[   472] = 11'd28;    
		mem[   473] = 11'd108;    
		mem[   474] = 11'd83;    
		mem[   475] = 11'd27;    
		mem[   476] = 11'd109;    
		mem[   477] = 11'd82;    
		mem[   478] = 11'd28;    
		mem[   479] = 11'd108;    
		mem[   480] = 11'd83;    
		mem[   481] = 11'd28;    
		mem[   482] = 11'd108;    
		mem[   483] = 11'd82;    
		mem[   484] = 11'd28;    
		mem[   485] = 11'd108;    
		mem[   486] = 11'd83;    
		mem[   487] = 11'd28;    
		mem[   488] = 11'd108;    
		mem[   489] = 11'd82;    
		mem[   490] = 11'd27;    
		mem[   491] = 11'd109;    
		mem[   492] = 11'd83;    
		mem[   493] = 11'd27;    
		mem[   494] = 11'd109;    
		mem[   495] = 11'd82;    
		mem[   496] = 11'd28;    
		mem[   497] = 11'd108;    
		mem[   498] = 11'd83;    
		mem[   499] = 11'd27;    
		mem[   500] = 11'd108;    
		mem[   501] = 11'd83;    
		mem[   502] = 11'd28;    
		mem[   503] = 11'd108;    
		mem[   504] = 11'd83;    
		mem[   505] = 11'd41;    
		mem[   506] = 11'd36;    
		mem[   507] = 11'd47;    
		mem[   508] = 11'd38;    
		mem[   509] = 11'd32;    
		mem[   510] = 11'd36;    
		mem[   511] = 11'd49;    
		mem[   512] = 11'd31;    
		mem[   513] = 11'd39;    
		mem[   514] = 11'd82;    
		mem[   515] = 11'd40;    
		mem[   516] = 11'd33;    
		mem[   517] = 11'd36;    
		mem[   518] = 11'd49;    
		mem[   519] = 11'd31;    
		mem[   520] = 11'd40;    
		mem[   521] = 11'd35;    
		mem[   522] = 11'd48;    
		mem[   523] = 11'd39;    
		mem[   524] = 11'd33;    
		mem[   525] = 11'd37;    
		mem[   526] = 11'd48;    
		mem[   527] = 11'd31;    
		mem[   528] = 11'd40;    
		mem[   529] = 11'd35;    
		mem[   530] = 11'd48;    
		mem[   531] = 11'd39;    
		mem[   532] = 11'd33;    
		mem[   533] = 11'd37;    
		mem[   534] = 11'd47;    
		mem[   535] = 11'd32;    
		mem[   536] = 11'd40;    
		mem[   537] = 11'd36;    
		mem[   538] = 11'd46;    
		mem[   539] = 11'd40;    
		mem[   540] = 11'd33;    
		mem[   541] = 11'd37;    
		mem[   542] = 11'd74;    
		mem[   543] = 11'd40;    
		mem[   544] = 11'd150;    
		mem[   545] = 11'd117;    
		mem[   546] = 11'd39;    
		mem[   547] = 11'd154;    
		mem[   548] = 11'd118;    
		mem[   549] = 11'd39;    
		mem[   550] = 11'd155;    
		mem[   551] = 11'd117;    
		mem[   552] = 11'd39;    
		mem[   553] = 11'd154;    
		mem[   554] = 11'd118;    
		mem[   555] = 11'd39;    
		mem[   556] = 11'd107;    
		mem[   557] = 11'd19;    
		mem[   558] = 11'd19;    
		mem[   559] = 11'd19;    
		mem[   560] = 11'd18;    
		mem[   561] = 11'd20;    
		mem[   562] = 11'd21;    
		mem[   563] = 11'd20;    
		mem[   564] = 11'd19;    
		mem[   565] = 11'd18;    
		mem[   566] = 11'd21;    
		mem[   567] = 11'd18;    
		mem[   568] = 11'd19;    
		mem[   569] = 11'd19;    
		mem[   570] = 11'd20;    
		mem[   571] = 11'd21;    
		mem[   572] = 11'd20;    
		mem[   573] = 11'd19;    
		mem[   574] = 11'd18;    
		mem[   575] = 11'd19;    
		mem[   576] = 11'd19;    
		mem[   577] = 11'd19;    
		mem[   578] = 11'd21;    
		mem[   579] = 11'd19;    
		mem[   580] = 11'd19;    
		mem[   581] = 11'd19;    
		mem[   582] = 11'd20;    
		mem[   583] = 11'd19;    
		mem[   584] = 11'd18;    
		mem[   585] = 11'd20;    
		mem[   586] = 11'd19;    
		mem[   587] = 11'd20;    
		mem[   588] = 11'd20;    
		mem[   589] = 11'd20;    
		mem[   590] = 11'd19;    
		mem[   591] = 11'd18;    
		mem[   592] = 11'd19;    
		mem[   593] = 11'd19;    
		mem[   594] = 11'd20;    
		mem[   595] = 11'd20;    
		mem[   596] = 11'd20;    
		mem[   597] = 11'd18;    
		mem[   598] = 11'd20;    
		mem[   599] = 11'd19;    
		mem[   600] = 11'd19;    
		mem[   601] = 11'd19;    
		mem[   602] = 11'd20;    
		mem[   603] = 11'd20;    
		mem[   604] = 11'd19;    
		mem[   605] = 11'd20;    
		mem[   606] = 11'd19;    
		mem[   607] = 11'd18;    
		mem[   608] = 11'd19;    
		mem[   609] = 11'd20;    
		mem[   610] = 11'd20;    
		mem[   611] = 11'd20;    
		mem[   612] = 11'd19;    
		mem[   613] = 11'd18;    
		mem[   614] = 11'd20;    
		mem[   615] = 11'd19;    
		mem[   616] = 11'd19;    
		mem[   617] = 11'd19;    
		mem[   618] = 11'd20;    
		mem[   619] = 11'd20;    
		mem[   620] = 11'd19;    
		mem[   621] = 11'd20;    
		mem[   622] = 11'd19;    
		mem[   623] = 11'd19;    
		mem[   624] = 11'd18;    
		mem[   625] = 11'd20;    
		mem[   626] = 11'd20;    
		mem[   627] = 11'd20;    
		mem[   628] = 11'd19;    
		mem[   629] = 11'd19;    
		mem[   630] = 11'd19;    
		mem[   631] = 11'd19;    
		mem[   632] = 11'd279;    
		mem[   633] = 11'd878;    
		mem[   634] = 11'd354;    
		mem[   635] = 11'd24;    
		mem[   636] = 11'd25;    
		mem[   637] = 11'd25;    
		mem[   638] = 11'd25;    
		mem[   639] = 11'd26;    
		mem[   640] = 11'd25;    
		mem[   641] = 11'd26;    
		mem[   642] = 11'd25;    
		mem[   643] = 11'd26;    
		mem[   644] = 11'd26;    
		mem[   645] = 11'd26;    
		mem[   646] = 11'd25;    
		mem[   647] = 11'd26;    
		mem[   648] = 11'd26;    
		mem[   649] = 11'd26;    
		mem[   650] = 11'd26;    
		mem[   651] = 11'd25;    
		mem[   652] = 11'd26;    
		mem[   653] = 11'd26;    
		mem[   654] = 11'd26;    
		mem[   655] = 11'd26;    
		mem[   656] = 11'd26;    
		mem[   657] = 11'd26;    
		mem[   658] = 11'd25;    
		mem[   659] = 11'd26;    
		mem[   660] = 11'd26;    
		mem[   661] = 11'd26;    
		mem[   662] = 11'd26;    
		mem[   663] = 11'd25;    
		mem[   664] = 11'd26;    
		mem[   665] = 11'd26;    
		mem[   666] = 11'd26;    
		mem[   667] = 11'd26;    
		mem[   668] = 11'd26;    
		mem[   669] = 11'd26;    
		mem[   670] = 11'd25;    
		mem[   671] = 11'd26;    
		mem[   672] = 11'd26;    
		mem[   673] = 11'd26;    
		mem[   674] = 11'd26;    
		mem[   675] = 11'd26;    
		mem[   676] = 11'd25;    
		mem[   677] = 11'd26;    
		mem[   678] = 11'd26;    
		mem[   679] = 11'd26;    
		mem[   680] = 11'd26;    
		mem[   681] = 11'd25;    
		mem[   682] = 11'd26;    
		mem[   683] = 11'd26;    
		mem[   684] = 11'd26;    
		mem[   685] = 11'd26;    
		mem[   686] = 11'd26;    
		mem[   687] = 11'd25;    
		mem[   688] = 11'd26;    
		mem[   689] = 11'd211;    
		mem[   690] = 11'd1272;    
		mem[   691] = 11'd28;    
		mem[   692] = 11'd30;    
		mem[   693] = 11'd69;    
		mem[   694] = 11'd27;    
		mem[   695] = 11'd66;    
		mem[   696] = 11'd21;    
		mem[   697] = 11'd18;    
		mem[   698] = 11'd14;    
		mem[   699] = 11'd34;    
		mem[   700] = 11'd36;    
		mem[   701] = 11'd25;    
		mem[   702] = 11'd30;    
		mem[   703] = 11'd35;    
		mem[   704] = 11'd31;    
		mem[   705] = 11'd23;    
		mem[   706] = 11'd37;    
		mem[   707] = 11'd32;    
		mem[   708] = 11'd24;    
		mem[   709] = 11'd37;    
		mem[   710] = 11'd29;    
		mem[   711] = 11'd29;    
		mem[   712] = 11'd26;    
		mem[   713] = 11'd39;    
		mem[   714] = 11'd29;    
		mem[   715] = 11'd24;    
		mem[   716] = 11'd39;    
		mem[   717] = 11'd26;    
		mem[   718] = 11'd30;    
		mem[   719] = 11'd30;    
		mem[   720] = 11'd37;    
		mem[   721] = 11'd27;    
		mem[   722] = 11'd26;    
		mem[   723] = 11'd38;    
		mem[   724] = 11'd22;    
		mem[   725] = 11'd33;    
		mem[   726] = 11'd33;    
		mem[   727] = 11'd35;    
		mem[   728] = 11'd25;    
		mem[   729] = 11'd31;    
		mem[   730] = 11'd34;    
		mem[   731] = 11'd31;    
		mem[   732] = 11'd25;    
		mem[   733] = 11'd36;    
		mem[   734] = 11'd31;    
		mem[   735] = 11'd25;    
		mem[   736] = 11'd36;    
		mem[   737] = 11'd54;    
		mem[   738] = 11'd104;    
		mem[   739] = 11'd79;    
		mem[   740] = 11'd29;    
		mem[   741] = 11'd103;    
		mem[   742] = 11'd78;    
		mem[   743] = 11'd26;    
		mem[   744] = 11'd103;    
		mem[   745] = 11'd77;    
		mem[   746] = 11'd26;    
		mem[   747] = 11'd100;    
		mem[   748] = 11'd77;    
		mem[   749] = 11'd27;    
		mem[   750] = 11'd102;    
		mem[   751] = 11'd77;    
		mem[   752] = 11'd27;    
		mem[   753] = 11'd102;    
		mem[   754] = 11'd78;    
		mem[   755] = 11'd29;    
		mem[   756] = 11'd100;    
		mem[   757] = 11'd84;    
		mem[   758] = 11'd18;    
		mem[   759] = 11'd19;    
		mem[   760] = 11'd17;    
		mem[   761] = 11'd19;    
		mem[   762] = 11'd19;    
		mem[   763] = 11'd22;    
		mem[   764] = 11'd22;    
		mem[   765] = 11'd36;    
		mem[   766] = 11'd18;    
		mem[   767] = 11'd17;    
		mem[   768] = 11'd39;    
		mem[   769] = 11'd24;    
		mem[   770] = 11'd19;    
		mem[   771] = 11'd17;    
		mem[   772] = 11'd40;    
		mem[   773] = 11'd15;    
		mem[   774] = 11'd39;    
		mem[   775] = 11'd21;    
		mem[   776] = 11'd22;    
		mem[   777] = 11'd20;    
		mem[   778] = 11'd18;    
		mem[   779] = 11'd18;    
		mem[   780] = 11'd16;    
		mem[   781] = 11'd41;    
		mem[   782] = 11'd22;    
		mem[   783] = 11'd20;    
		mem[   784] = 11'd18;    
		mem[   785] = 11'd12;    
		mem[   786] = 11'd27;    
		mem[   787] = 11'd16;    
		mem[   788] = 11'd38;    
		mem[   789] = 11'd21;    
		mem[   790] = 11'd22;    
		mem[   791] = 11'd20;    
		mem[   792] = 11'd19;    
		mem[   793] = 11'd18;    
		mem[   794] = 11'd16;    
		mem[   795] = 11'd40;    
		mem[   796] = 11'd22;    
		mem[   797] = 11'd20;    
		mem[   798] = 11'd18;    
		mem[   799] = 11'd15;    
		mem[   800] = 11'd25;    
		mem[   801] = 11'd16;    
		mem[   802] = 11'd18;    
		mem[   803] = 11'd20;    
		mem[   804] = 11'd21;    
		mem[   805] = 11'd21;    
		mem[   806] = 11'd20;    
		mem[   807] = 11'd19;    
		mem[   808] = 11'd18;    
		mem[   809] = 11'd17;    
		mem[   810] = 11'd18;    
		mem[   811] = 11'd21;    
		mem[   812] = 11'd22;    
		mem[   813] = 11'd20;    
		mem[   814] = 11'd18;    
		mem[   815] = 11'd16;    
		mem[   816] = 11'd24;    
		mem[   817] = 11'd16;    
		mem[   818] = 11'd18;    
		mem[   819] = 11'd20;    
		mem[   820] = 11'd21;    
		mem[   821] = 11'd21;    
		mem[   822] = 11'd20;    
		mem[   823] = 11'd19;    
		mem[   824] = 11'd18;    
		mem[   825] = 11'd18;    
		mem[   826] = 11'd25;    
		mem[   827] = 11'd29;    
		mem[   828] = 11'd29;    
		mem[   829] = 11'd23;    
		mem[   830] = 11'd25;    
		mem[   831] = 11'd25;    
		mem[   832] = 11'd24;    
		mem[   833] = 11'd28;    
		mem[   834] = 11'd28;    
		mem[   835] = 11'd28;    
		mem[   836] = 11'd24;    
		mem[   837] = 11'd22;    
		mem[   838] = 11'd24;    
		mem[   839] = 11'd30;    
		mem[   840] = 11'd28;    
		mem[   841] = 11'd24;    
		mem[   842] = 11'd25;    
		mem[   843] = 11'd25;    
		mem[   844] = 11'd24;    
		mem[   845] = 11'd27;    
		mem[   846] = 11'd29;    
		mem[   847] = 11'd27;    
		mem[   848] = 11'd24;    
		mem[   849] = 11'd23;    
		mem[   850] = 11'd25;    
		mem[   851] = 11'd29;    
		mem[   852] = 11'd28;    
		mem[   853] = 11'd24;    
		mem[   854] = 11'd24;    
		mem[   855] = 11'd26;    
		mem[   856] = 11'd24;    
		mem[   857] = 11'd27;    
		mem[   858] = 11'd28;    
		mem[   859] = 11'd27;    
		mem[   860] = 11'd25;    
		mem[   861] = 11'd23;    
		mem[   862] = 11'd25;    
		mem[   863] = 11'd29;    
		mem[   864] = 11'd27;    
		mem[   865] = 11'd25;    
		mem[   866] = 11'd24;    
		mem[   867] = 11'd26;    
		mem[   868] = 11'd24;    
		mem[   869] = 11'd27;    
		mem[   870] = 11'd28;    
		mem[   871] = 11'd26;    
		mem[   872] = 11'd25;    
		mem[   873] = 11'd25;    
		mem[   874] = 11'd24;    
		mem[   875] = 11'd28;    
		mem[   876] = 11'd27;    
		mem[   877] = 11'd25;    
		mem[   878] = 11'd25;    
		mem[   879] = 11'd26;    
		mem[   880] = 11'd24;    
		mem[   881] = 11'd27;    
		mem[   882] = 11'd213;    
		mem[   883] = 11'd47;    
		mem[   884] = 11'd156;    
		mem[   885] = 11'd116;    
		mem[   886] = 11'd39;    
		mem[   887] = 11'd154;    
		mem[   888] = 11'd112;    
		mem[   889] = 11'd40;    
		mem[   890] = 11'd152;    
		mem[   891] = 11'd116;    
		mem[   892] = 11'd42;    
		mem[   893] = 11'd154;    
		mem[   894] = 11'd115;    
		mem[   895] = 11'd39;    
		mem[   896] = 11'd154;    
		mem[   897] = 11'd120;    
		mem[   898] = 11'd38;    
		mem[   899] = 11'd154;    
		mem[   900] = 11'd125;    
		mem[   901] = 11'd39;    
		mem[   902] = 11'd823;    
		mem[   903] = 11'd29;    
		mem[   904] = 11'd30;    
		mem[   905] = 11'd30;    
		mem[   906] = 11'd30;    
		mem[   907] = 11'd30;    
		mem[   908] = 11'd31;    
		mem[   909] = 11'd30;    
		mem[   910] = 11'd31;    
		mem[   911] = 11'd30;    
		mem[   912] = 11'd31;    
		mem[   913] = 11'd30;    
		mem[   914] = 11'd31;    
		mem[   915] = 11'd31;    
		mem[   916] = 11'd31;    
		mem[   917] = 11'd30;    
		mem[   918] = 11'd31;    
		mem[   919] = 11'd30;    
		mem[   920] = 11'd31;    
		mem[   921] = 11'd31;    
		mem[   922] = 11'd30;    
		mem[   923] = 11'd31;    
		mem[   924] = 11'd31;    
		mem[   925] = 11'd30;    
		mem[   926] = 11'd31;    
		mem[   927] = 11'd31;    
		mem[   928] = 11'd30;    
		mem[   929] = 11'd31;    
		mem[   930] = 11'd31;    
		mem[   931] = 11'd30;    
		mem[   932] = 11'd31;    
		mem[   933] = 11'd31;    
		mem[   934] = 11'd30;    
		mem[   935] = 11'd31;    
		mem[   936] = 11'd31;    
		mem[   937] = 11'd30;    
		mem[   938] = 11'd31;    
		mem[   939] = 11'd31;    
		mem[   940] = 11'd30;    
		mem[   941] = 11'd31;    
		mem[   942] = 11'd30;    
		mem[   943] = 11'd31;    
		mem[   944] = 11'd31;    
		mem[   945] = 11'd30;    
		mem[   946] = 11'd31;    
		mem[   947] = 11'd31;    
		mem[   948] = 11'd30;    
		mem[   949] = 11'd31;    
		mem[   950] = 11'd31;    
		mem[   951] = 11'd30;    
		mem[   952] = 11'd31;    
		mem[   953] = 11'd31;    
		mem[   954] = 11'd30;    
		mem[   955] = 11'd31;    
		mem[   956] = 11'd30;    
		mem[   957] = 11'd31;    
		mem[   958] = 11'd31;    
		mem[   959] = 11'd30;    
		mem[   960] = 11'd31;    
		mem[   961] = 11'd31;    
		mem[   962] = 11'd30;    
		mem[   963] = 11'd31;    
		mem[   964] = 11'd31;    
		mem[   965] = 11'd30;    
		mem[   966] = 11'd31;    
		mem[   967] = 11'd30;    
		mem[   968] = 11'd31;    
		mem[   969] = 11'd31;    
		mem[   970] = 11'd30;    
		mem[   971] = 11'd31;    
		mem[   972] = 11'd31;    
		mem[   973] = 11'd30;    
		mem[   974] = 11'd31;    
		mem[   975] = 11'd31;    
		mem[   976] = 11'd30;    
		mem[   977] = 11'd31;    
		mem[   978] = 11'd30;    
		mem[   979] = 11'd31;    
		mem[   980] = 11'd31;    
		mem[   981] = 11'd30;    
		mem[   982] = 11'd31;    
		mem[   983] = 11'd31;    
		mem[   984] = 11'd30;    
		mem[   985] = 11'd31;    
		mem[   986] = 11'd31;    
		mem[   987] = 11'd30;    
		mem[   988] = 11'd31;    
		mem[   989] = 11'd31;    
		mem[   990] = 11'd30;    
		mem[   991] = 11'd31;    
		mem[   992] = 11'd30;    
		mem[   993] = 11'd31;    
		mem[   994] = 11'd31;    
		mem[   995] = 11'd30;    
		mem[   996] = 11'd31;    
		mem[   997] = 11'd70;    
		mem[   998] = 11'd27;    
		mem[   999] = 11'd102;    
		mem[  1000] = 11'd78;    
		mem[  1001] = 11'd27;    
		mem[  1002] = 11'd101;    
		mem[  1003] = 11'd78;    
		mem[  1004] = 11'd27;    
		mem[  1005] = 11'd102;    
		mem[  1006] = 11'd78;    
		mem[  1007] = 11'd26;    
		mem[  1008] = 11'd102;    
		mem[  1009] = 11'd79;    
		mem[  1010] = 11'd26;    
		mem[  1011] = 11'd102;    
		mem[  1012] = 11'd78;    
		mem[  1013] = 11'd26;    
		mem[  1014] = 11'd102;    
		mem[  1015] = 11'd78;    
		mem[  1016] = 11'd26;    
		mem[  1017] = 11'd103;    
		mem[  1018] = 11'd78;    
		mem[  1019] = 11'd26;    
		mem[  1020] = 11'd103;    
		mem[  1021] = 11'd77;    
		mem[  1022] = 11'd27;    
		mem[  1023] = 11'd102;    
		mem[  1024] = 11'd78;    
		mem[  1025] = 11'd26;    
		mem[  1026] = 11'd102;    
		mem[  1027] = 11'd78;    
		mem[  1028] = 11'd27;    
		mem[  1029] = 11'd102;    
		mem[  1030] = 11'd78;    
		mem[  1031] = 11'd26;    
		mem[  1032] = 11'd102;    
		mem[  1033] = 11'd78;    
		mem[  1034] = 11'd26;    
		mem[  1035] = 11'd103;    
		mem[  1036] = 11'd78;    
		mem[  1037] = 11'd26;    
		mem[  1038] = 11'd103;    
		mem[  1039] = 11'd107;    
		mem[  1040] = 11'd41;    
		mem[  1041] = 11'd37;    
		mem[  1042] = 11'd50;    
		mem[  1043] = 11'd41;    
		mem[  1044] = 11'd35;    
		mem[  1045] = 11'd37;    
		mem[  1046] = 11'd52;    
		mem[  1047] = 11'd33;    
		mem[  1048] = 11'd42;    
		mem[  1049] = 11'd34;    
		mem[  1050] = 11'd53;    
		mem[  1051] = 11'd41;    
		mem[  1052] = 11'd35;    
		mem[  1053] = 11'd38;    
		mem[  1054] = 11'd52;    
		mem[  1055] = 11'd33;    
		mem[  1056] = 11'd42;    
		mem[  1057] = 11'd36;    
		mem[  1058] = 11'd50;    
		mem[  1059] = 11'd42;    
		mem[  1060] = 11'd35;    
		mem[  1061] = 11'd39;    
		mem[  1062] = 11'd50;    
		mem[  1063] = 11'd34;    
		mem[  1064] = 11'd42;    
		mem[  1065] = 11'd37;    
		mem[  1066] = 11'd49;    
		mem[  1067] = 11'd41;    
		mem[  1068] = 11'd36;    
		mem[  1069] = 11'd39;    
		mem[  1070] = 11'd49;    
		mem[  1071] = 11'd35;    
		mem[  1072] = 11'd41;    
		mem[  1073] = 11'd38;    
		mem[  1074] = 11'd117;    
		mem[  1075] = 11'd122;    
		mem[  1076] = 11'd42;    
		mem[  1077] = 11'd162;    
		mem[  1078] = 11'd124;    
		mem[  1079] = 11'd41;    
		mem[  1080] = 11'd163;    
		mem[  1081] = 11'd124;    
		mem[  1082] = 11'd42;    
		mem[  1083] = 11'd161;    
		mem[  1084] = 11'd124;    
		mem[  1085] = 11'd42;    
		mem[  1086] = 11'd163;    
		mem[  1087] = 11'd53;    
		mem[  1088] = 11'd22;    
		mem[  1089] = 11'd21;    
		mem[  1090] = 11'd20;    
		mem[  1091] = 11'd19;    
		mem[  1092] = 11'd23;    
		mem[  1093] = 11'd19;    
		mem[  1094] = 11'd20;    
		mem[  1095] = 11'd21;    
		mem[  1096] = 11'd21;    
		mem[  1097] = 11'd21;    
		mem[  1098] = 11'd21;    
		mem[  1099] = 11'd20;    
		mem[  1100] = 11'd20;    
		mem[  1101] = 11'd20;    
		mem[  1102] = 11'd20;    
		mem[  1103] = 11'd21;    
		mem[  1104] = 11'd22;    
		mem[  1105] = 11'd20;    
		mem[  1106] = 11'd20;    
		mem[  1107] = 11'd19;    
		mem[  1108] = 11'd23;    
		mem[  1109] = 11'd19;    
		mem[  1110] = 11'd20;    
		mem[  1111] = 11'd21;    
		mem[  1112] = 11'd21;    
		mem[  1113] = 11'd21;    
		mem[  1114] = 11'd21;    
		mem[  1115] = 11'd20;    
		mem[  1116] = 11'd20;    
		mem[  1117] = 11'd19;    
		mem[  1118] = 11'd20;    
		mem[  1119] = 11'd22;    
		mem[  1120] = 11'd21;    
		mem[  1121] = 11'd21;    
		mem[  1122] = 11'd20;    
		mem[  1123] = 11'd19;    
		mem[  1124] = 11'd22;    
		mem[  1125] = 11'd19;    
		mem[  1126] = 11'd21;    
		mem[  1127] = 11'd20;    
		mem[  1128] = 11'd21;    
		mem[  1129] = 11'd21;    
		mem[  1130] = 11'd21;    
		mem[  1131] = 11'd20;    
		mem[  1132] = 11'd20;    
		mem[  1133] = 11'd20;    
		mem[  1134] = 11'd20;    
		mem[  1135] = 11'd21;    
		mem[  1136] = 11'd22;    
		mem[  1137] = 11'd20;    
		mem[  1138] = 11'd20;    
		mem[  1139] = 11'd20;    
		mem[  1140] = 11'd22;    
		mem[  1141] = 11'd19;    
		mem[  1142] = 11'd20;    
		mem[  1143] = 11'd21;    
		mem[  1144] = 11'd21;    
		mem[  1145] = 11'd21;    
		mem[  1146] = 11'd20;    
		mem[  1147] = 11'd21;    
		mem[  1148] = 11'd20;    
		mem[  1149] = 11'd20;    
		mem[  1150] = 11'd20;    
		mem[  1151] = 11'd21;    
		mem[  1152] = 11'd21;    
		mem[  1153] = 11'd21;    
		mem[  1154] = 11'd20;    
		mem[  1155] = 11'd20;    
		mem[  1156] = 11'd21;    
		mem[  1157] = 11'd20;    
		mem[  1158] = 11'd282;    
		mem[  1159] = 11'd44;    
		mem[  1160] = 11'd174;    
		mem[  1161] = 11'd112;    
		mem[  1162] = 11'd42;    
		mem[  1163] = 11'd334;    
		mem[  1164] = 11'd527;    
		mem[  1165] = 11'd26;    
		mem[  1166] = 11'd26;    
		mem[  1167] = 11'd27;    
		mem[  1168] = 11'd27;    
		mem[  1169] = 11'd27;    
		mem[  1170] = 11'd27;    
		mem[  1171] = 11'd27;    
		mem[  1172] = 11'd27;    
		mem[  1173] = 11'd27;    
		mem[  1174] = 11'd27;    
		mem[  1175] = 11'd27;    
		mem[  1176] = 11'd28;    
		mem[  1177] = 11'd27;    
		mem[  1178] = 11'd27;    
		mem[  1179] = 11'd28;    
		mem[  1180] = 11'd27;    
		mem[  1181] = 11'd27;    
		mem[  1182] = 11'd28;    
		mem[  1183] = 11'd27;    
		mem[  1184] = 11'd27;    
		mem[  1185] = 11'd28;    
		mem[  1186] = 11'd27;    
		mem[  1187] = 11'd27;    
		mem[  1188] = 11'd28;    
		mem[  1189] = 11'd27;    
		mem[  1190] = 11'd28;    
		mem[  1191] = 11'd27;    
		mem[  1192] = 11'd27;    
		mem[  1193] = 11'd27;    
		mem[  1194] = 11'd28;    
		mem[  1195] = 11'd27;    
		mem[  1196] = 11'd27;    
		mem[  1197] = 11'd28;    
		mem[  1198] = 11'd27;    
		mem[  1199] = 11'd27;    
		mem[  1200] = 11'd28;    
		mem[  1201] = 11'd27;    
		mem[  1202] = 11'd28;    
		mem[  1203] = 11'd27;    
		mem[  1204] = 11'd27;    
		mem[  1205] = 11'd27;    
		mem[  1206] = 11'd28;    
		mem[  1207] = 11'd27;    
		mem[  1208] = 11'd27;    
		mem[  1209] = 11'd28;    
		mem[  1210] = 11'd27;    
		mem[  1211] = 11'd27;    
		mem[  1212] = 11'd28;    
		mem[  1213] = 11'd27;    
		mem[  1214] = 11'd27;    
		mem[  1215] = 11'd28;    
		mem[  1216] = 11'd1484;    
		mem[  1217] = 11'd69;    
		mem[  1218] = 11'd31;    
		mem[  1219] = 11'd27;    
		mem[  1220] = 11'd43;    
		mem[  1221] = 11'd29;    
		mem[  1222] = 11'd25;    
		mem[  1223] = 11'd44;    
		mem[  1224] = 11'd25;    
		mem[  1225] = 11'd32;    
		mem[  1226] = 11'd32;    
		mem[  1227] = 11'd41;    
		mem[  1228] = 11'd26;    
		mem[  1229] = 11'd29;    
		mem[  1230] = 11'd40;    
		mem[  1231] = 11'd21;    
		mem[  1232] = 11'd8;    
		mem[  1233] = 11'd29;    
		mem[  1234] = 11'd37;    
		mem[  1235] = 11'd36;    
		mem[  1236] = 11'd25;    
		mem[  1237] = 11'd36;    
		mem[  1238] = 11'd34;    
		mem[  1239] = 11'd32;    
		mem[  1240] = 11'd27;    
		mem[  1241] = 11'd39;    
		mem[  1242] = 11'd33;    
		mem[  1243] = 11'd25;    
		mem[  1244] = 11'd41;    
		mem[  1245] = 11'd28;    
		mem[  1246] = 11'd32;    
		mem[  1247] = 11'd30;    
		mem[  1248] = 11'd40;    
		mem[  1249] = 11'd29;    
		mem[  1250] = 11'd27;    
		mem[  1251] = 11'd42;    
		mem[  1252] = 11'd24;    
		mem[  1253] = 11'd34;    
		mem[  1254] = 11'd34;    
		mem[  1255] = 11'd38;    
		mem[  1256] = 11'd28;    
		mem[  1257] = 11'd31;    
		mem[  1258] = 11'd37;    
		mem[  1259] = 11'd16;    
		mem[  1260] = 11'd17;    
		mem[  1261] = 11'd25;    
		mem[  1262] = 11'd79;    
		mem[  1263] = 11'd91;    
		mem[  1264] = 11'd28;    
		mem[  1265] = 11'd112;    
		mem[  1266] = 11'd80;    
		mem[  1267] = 11'd31;    
		mem[  1268] = 11'd108;    
		mem[  1269] = 11'd82;    
		mem[  1270] = 11'd28;    
		mem[  1271] = 11'd105;    
		mem[  1272] = 11'd82;    
		mem[  1273] = 11'd30;    
		mem[  1274] = 11'd106;    
		mem[  1275] = 11'd82;    
		mem[  1276] = 11'd28;    
		mem[  1277] = 11'd108;    
		mem[  1278] = 11'd82;    
		mem[  1279] = 11'd29;    
		mem[  1280] = 11'd108;    
		mem[  1281] = 11'd90;    
		mem[  1282] = 11'd20;    
		mem[  1283] = 11'd20;    
		mem[  1284] = 11'd17;    
		mem[  1285] = 11'd20;    
		mem[  1286] = 11'd21;    
		mem[  1287] = 11'd23;    
		mem[  1288] = 11'd23;    
		mem[  1289] = 11'd21;    
		mem[  1290] = 11'd18;    
		mem[  1291] = 11'd18;    
		mem[  1292] = 11'd18;    
		mem[  1293] = 11'd44;    
		mem[  1294] = 11'd23;    
		mem[  1295] = 11'd20;    
		mem[  1296] = 11'd18;    
		mem[  1297] = 11'd41;    
		mem[  1298] = 11'd18;    
		mem[  1299] = 11'd41;    
		mem[  1300] = 11'd24;    
		mem[  1301] = 11'd22;    
		mem[  1302] = 11'd21;    
		mem[  1303] = 11'd19;    
		mem[  1304] = 11'd18;    
		mem[  1305] = 11'd18;    
		mem[  1306] = 11'd45;    
		mem[  1307] = 11'd23;    
		mem[  1308] = 11'd19;    
		mem[  1309] = 11'd18;    
		mem[  1310] = 11'd42;    
		mem[  1311] = 11'd18;    
		mem[  1312] = 11'd20;    
		mem[  1313] = 11'd21;    
		mem[  1314] = 11'd23;    
		mem[  1315] = 11'd23;    
		mem[  1316] = 11'd21;    
		mem[  1317] = 11'd19;    
		mem[  1318] = 11'd18;    
		mem[  1319] = 11'd19;    
		mem[  1320] = 11'd43;    
		mem[  1321] = 11'd23;    
		mem[  1322] = 11'd20;    
		mem[  1323] = 11'd18;    
		mem[  1324] = 11'd41;    
		mem[  1325] = 11'd19;    
		mem[  1326] = 11'd20;    
		mem[  1327] = 11'd21;    
		mem[  1328] = 11'd23;    
		mem[  1329] = 11'd22;    
		mem[  1330] = 11'd21;    
		mem[  1331] = 11'd19;    
		mem[  1332] = 11'd19;    
		mem[  1333] = 11'd19;    
		mem[  1334] = 11'd19;    
		mem[  1335] = 11'd24;    
		mem[  1336] = 11'd23;    
		mem[  1337] = 11'd20;    
		mem[  1338] = 11'd18;    
		mem[  1339] = 11'd17;    
		mem[  1340] = 11'd24;    
		mem[  1341] = 11'd19;    
		mem[  1342] = 11'd20;    
		mem[  1343] = 11'd21;    
		mem[  1344] = 11'd23;    
		mem[  1345] = 11'd26;    
		mem[  1346] = 11'd27;    
		mem[  1347] = 11'd25;    
		mem[  1348] = 11'd24;    
		mem[  1349] = 11'd29;    
		mem[  1350] = 11'd32;    
		mem[  1351] = 11'd26;    
		mem[  1352] = 11'd23;    
		mem[  1353] = 11'd31;    
		mem[  1354] = 11'd23;    
		mem[  1355] = 11'd28;    
		mem[  1356] = 11'd29;    
		mem[  1357] = 11'd30;    
		mem[  1358] = 11'd27;    
		mem[  1359] = 11'd26;    
		mem[  1360] = 11'd24;    
		mem[  1361] = 11'd29;    
		mem[  1362] = 11'd31;    
		mem[  1363] = 11'd26;    
		mem[  1364] = 11'd24;    
		mem[  1365] = 11'd30;    
		mem[  1366] = 11'd24;    
		mem[  1367] = 11'd28;    
		mem[  1368] = 11'd29;    
		mem[  1369] = 11'd30;    
		mem[  1370] = 11'd27;    
		mem[  1371] = 11'd25;    
		mem[  1372] = 11'd25;    
		mem[  1373] = 11'd28;    
		mem[  1374] = 11'd31;    
		mem[  1375] = 11'd27;    
		mem[  1376] = 11'd24;    
		mem[  1377] = 11'd30;    
		mem[  1378] = 11'd24;    
		mem[  1379] = 11'd27;    
		mem[  1380] = 11'd30;    
		mem[  1381] = 11'd29;    
		mem[  1382] = 11'd27;    
		mem[  1383] = 11'd26;    
		mem[  1384] = 11'd24;    
		mem[  1385] = 11'd29;    
		mem[  1386] = 11'd30;    
		mem[  1387] = 11'd27;    
		mem[  1388] = 11'd25;    
		mem[  1389] = 11'd30;    
		mem[  1390] = 11'd24;    
		mem[  1391] = 11'd28;    
		mem[  1392] = 11'd28;    
		mem[  1393] = 11'd30;    
		mem[  1394] = 11'd27;    
		mem[  1395] = 11'd26;    
		mem[  1396] = 11'd25;    
		mem[  1397] = 11'd28;    
		mem[  1398] = 11'd83;    
		mem[  1399] = 11'd48;    
		mem[  1400] = 11'd141;    
		mem[  1401] = 11'd118;    
		mem[  1402] = 11'd50;    
		mem[  1403] = 11'd154;    
		mem[  1404] = 11'd132;    
		mem[  1405] = 11'd42;    
		mem[  1406] = 11'd162;    
		mem[  1407] = 11'd124;    
		mem[  1408] = 11'd42;    
		mem[  1409] = 11'd162;    
		mem[  1410] = 11'd124;    
		mem[  1411] = 11'd42;    
		mem[  1412] = 11'd164;    
		mem[  1413] = 11'd122;    
		mem[  1414] = 11'd44;    
		mem[  1415] = 11'd160;    
		mem[  1416] = 11'd124;    
		mem[  1417] = 11'd42;    
		mem[  1418] = 11'd130;    
		mem[  1419] = 11'd793;    
		mem[  1420] = 11'd35;    
		mem[  1421] = 11'd33;    
		mem[  1422] = 11'd34;    
		mem[  1423] = 11'd33;    
		mem[  1424] = 11'd32;    
		mem[  1425] = 11'd33;    
		mem[  1426] = 11'd33;    
		mem[  1427] = 11'd32;    
		mem[  1428] = 11'd33;    
		mem[  1429] = 11'd32;    
		mem[  1430] = 11'd33;    
		mem[  1431] = 11'd32;    
		mem[  1432] = 11'd33;    
		mem[  1433] = 11'd32;    
		mem[  1434] = 11'd33;    
		mem[  1435] = 11'd32;    
		mem[  1436] = 11'd32;    
		mem[  1437] = 11'd33;    
		mem[  1438] = 11'd32;    
		mem[  1439] = 11'd33;    
		mem[  1440] = 11'd32;    
		mem[  1441] = 11'd33;    
		mem[  1442] = 11'd32;    
		mem[  1443] = 11'd33;    
		mem[  1444] = 11'd32;    
		mem[  1445] = 11'd32;    
		mem[  1446] = 11'd33;    
		mem[  1447] = 11'd32;    
		mem[  1448] = 11'd33;    
		mem[  1449] = 11'd32;    
		mem[  1450] = 11'd33;    
		mem[  1451] = 11'd32;    
		mem[  1452] = 11'd33;    
		mem[  1453] = 11'd32;    
		mem[  1454] = 11'd33;    
		mem[  1455] = 11'd32;    
		mem[  1456] = 11'd33;    
		mem[  1457] = 11'd32;    
		mem[  1458] = 11'd32;    
		mem[  1459] = 11'd33;    
		mem[  1460] = 11'd32;    
		mem[  1461] = 11'd33;    
		mem[  1462] = 11'd32;    
		mem[  1463] = 11'd33;    
		mem[  1464] = 11'd32;    
		mem[  1465] = 11'd33;    
		mem[  1466] = 11'd32;    
		mem[  1467] = 11'd33;    
		mem[  1468] = 11'd32;    
		mem[  1469] = 11'd33;    
		mem[  1470] = 11'd32;    
		mem[  1471] = 11'd33;    
		mem[  1472] = 11'd32;    
		mem[  1473] = 11'd33;    
		mem[  1474] = 11'd32;    
		mem[  1475] = 11'd33;    
		mem[  1476] = 11'd32;    
		mem[  1477] = 11'd33;    
		mem[  1478] = 11'd32;    
		mem[  1479] = 11'd33;    
		mem[  1480] = 11'd32;    
		mem[  1481] = 11'd33;    
		mem[  1482] = 11'd32;    
		mem[  1483] = 11'd32;    
		mem[  1484] = 11'd33;    
		mem[  1485] = 11'd32;    
		mem[  1486] = 11'd33;    
		mem[  1487] = 11'd32;    
		mem[  1488] = 11'd33;    
		mem[  1489] = 11'd32;    
		mem[  1490] = 11'd33;    
		mem[  1491] = 11'd32;    
		mem[  1492] = 11'd33;    
		mem[  1493] = 11'd32;    
		mem[  1494] = 11'd33;    
		mem[  1495] = 11'd32;    
		mem[  1496] = 11'd33;    
		mem[  1497] = 11'd32;    
		mem[  1498] = 11'd33;    
		mem[  1499] = 11'd32;    
		mem[  1500] = 11'd33;    
		mem[  1501] = 11'd32;    
		mem[  1502] = 11'd33;    
		mem[  1503] = 11'd32;    
		mem[  1504] = 11'd33;    
		mem[  1505] = 11'd32;    
		mem[  1506] = 11'd33;    
		mem[  1507] = 11'd79;    
		mem[  1508] = 11'd28;    
		mem[  1509] = 11'd102;    
		mem[  1510] = 11'd82;    
		mem[  1511] = 11'd28;    
		mem[  1512] = 11'd107;    
		mem[  1513] = 11'd83;    
		mem[  1514] = 11'd28;    
		mem[  1515] = 11'd108;    
		mem[  1516] = 11'd83;    
		mem[  1517] = 11'd28;    
		mem[  1518] = 11'd108;    
		mem[  1519] = 11'd83;    
		mem[  1520] = 11'd28;    
		mem[  1521] = 11'd108;    
		mem[  1522] = 11'd82;    
		mem[  1523] = 11'd28;    
		mem[  1524] = 11'd109;    
		mem[  1525] = 11'd82;    
		mem[  1526] = 11'd28;    
		mem[  1527] = 11'd108;    
		mem[  1528] = 11'd83;    
		mem[  1529] = 11'd27;    
		mem[  1530] = 11'd109;    
		mem[  1531] = 11'd82;    
		mem[  1532] = 11'd28;    
		mem[  1533] = 11'd108;    
		mem[  1534] = 11'd83;    
		mem[  1535] = 11'd27;    
		mem[  1536] = 11'd109;    
		mem[  1537] = 11'd82;    
		mem[  1538] = 11'd27;    
		mem[  1539] = 11'd109;    
		mem[  1540] = 11'd82;    
		mem[  1541] = 11'd28;    
		mem[  1542] = 11'd108;    
		mem[  1543] = 11'd83;    
		mem[  1544] = 11'd30;    
		mem[  1545] = 11'd106;    
		mem[  1546] = 11'd83;    
		mem[  1547] = 11'd31;    
		mem[  1548] = 11'd76;    
		mem[  1549] = 11'd29;    
		mem[  1550] = 11'd31;    
		mem[  1551] = 11'd42;    
		mem[  1552] = 11'd34;    
		mem[  1553] = 11'd27;    
		mem[  1554] = 11'd45;    
		mem[  1555] = 11'd32;    
		mem[  1556] = 11'd26;    
		mem[  1557] = 11'd46;    
		mem[  1558] = 11'd24;    
		mem[  1559] = 11'd36;    
		mem[  1560] = 11'd39;    
		mem[  1561] = 11'd38;    
		mem[  1562] = 11'd27;    
		mem[  1563] = 11'd41;    
		mem[  1564] = 11'd31;    
		mem[  1565] = 11'd33;    
		mem[  1566] = 11'd34;    
		mem[  1567] = 11'd43;    
		mem[  1568] = 11'd28;    
		mem[  1569] = 11'd33;    
		mem[  1570] = 11'd39;    
		mem[  1571] = 11'd34;    
		mem[  1572] = 11'd28;    
		mem[  1573] = 11'd44;    
		mem[  1574] = 11'd32;    
		mem[  1575] = 11'd27;    
		mem[  1576] = 11'd45;    
		mem[  1577] = 11'd24;    
		mem[  1578] = 11'd37;    
		mem[  1579] = 11'd39;    
		mem[  1580] = 11'd37;    
		mem[  1581] = 11'd28;    
		mem[  1582] = 11'd41;    
		mem[  1583] = 11'd31;    
		mem[  1584] = 11'd33;    
		mem[  1585] = 11'd34;    
		mem[  1586] = 11'd42;    
		mem[  1587] = 11'd29;    
		mem[  1588] = 11'd33;    
		mem[  1589] = 11'd37;    
		mem[  1590] = 11'd32;    
		mem[  1591] = 11'd27;    
		mem[  1592] = 11'd37;    
		mem[  1593] = 11'd34;    
		mem[  1594] = 11'd27;    
		mem[  1595] = 11'd37;    
		mem[  1596] = 11'd31;    
		mem[  1597] = 11'd32;    
		mem[  1598] = 11'd29;    
		mem[  1599] = 11'd39;    
		mem[  1600] = 11'd31;    
		mem[  1601] = 11'd27;    
		mem[  1602] = 11'd39;    
		mem[  1603] = 11'd28;    
		mem[  1604] = 11'd33;    
		mem[  1605] = 11'd32;    
		mem[  1606] = 11'd38;    
		mem[  1607] = 11'd29;    
		mem[  1608] = 11'd30;    
		mem[  1609] = 11'd37;    
		mem[  1610] = 11'd30;    
		mem[  1611] = 11'd30;    
		mem[  1612] = 11'd35;    
		mem[  1613] = 11'd35;    
		mem[  1614] = 11'd28;    
		mem[  1615] = 11'd35;    
		mem[  1616] = 11'd34;    
		mem[  1617] = 11'd32;    
		mem[  1618] = 11'd28;    
		mem[  1619] = 11'd37;    
		mem[  1620] = 11'd33;    
		mem[  1621] = 11'd28;    
		mem[  1622] = 11'd36;    
		mem[  1623] = 11'd31;    
		mem[  1624] = 11'd32;    
		mem[  1625] = 11'd32;    
		mem[  1626] = 11'd36;    
		mem[  1627] = 11'd31;    
		mem[  1628] = 11'd30;    
		mem[  1629] = 11'd37;    
		mem[  1630] = 11'd28;    
		mem[  1631] = 11'd33;    
		mem[  1632] = 11'd33;    
		mem[  1633] = 11'd35;    
		mem[  1634] = 11'd28;    
		mem[  1635] = 11'd30;    
		mem[  1636] = 11'd33;    
		mem[  1637] = 11'd27;    
		mem[  1638] = 11'd32;    
		mem[  1639] = 11'd31;    
		mem[  1640] = 11'd33;    
		mem[  1641] = 11'd29;    
		mem[  1642] = 11'd29;    
		mem[  1643] = 11'd34;    
		mem[  1644] = 11'd28;    
		mem[  1645] = 11'd31;    
		mem[  1646] = 11'd30;    
		mem[  1647] = 11'd33;    
		mem[  1648] = 11'd30;    
		mem[  1649] = 11'd28;    
		mem[  1650] = 11'd34;    
		mem[  1651] = 11'd29;    
		mem[  1652] = 11'd30;    
		mem[  1653] = 11'd30;    
		mem[  1654] = 11'd33;    
		mem[  1655] = 11'd31;    
		mem[  1656] = 11'd28;    
		mem[  1657] = 11'd33;    
		mem[  1658] = 11'd30;    
		mem[  1659] = 11'd30;    
		mem[  1660] = 11'd30;    
		mem[  1661] = 11'd32;    
		mem[  1662] = 11'd31;    
		mem[  1663] = 11'd29;    
		mem[  1664] = 11'd32;    
		mem[  1665] = 11'd31;    
		mem[  1666] = 11'd30;    
		mem[  1667] = 11'd29;    
		mem[  1668] = 11'd32;    
		mem[  1669] = 11'd31;    
		mem[  1670] = 11'd30;    
		mem[  1671] = 11'd31;    
		mem[  1672] = 11'd31;    
		mem[  1673] = 11'd31;    
		mem[  1674] = 11'd29;    
		mem[  1675] = 11'd32;    
		mem[  1676] = 11'd31;    
		mem[  1677] = 11'd29;    
		mem[  1678] = 11'd31;    
		mem[  1679] = 11'd32;    
		mem[  1680] = 11'd30;    
		mem[  1681] = 11'd205;    
		mem[  1682] = 11'd31;    
		mem[  1683] = 11'd118;    
		mem[  1684] = 11'd838;    
		mem[  1685] = 11'd355;    
		mem[  1686] = 11'd34;    
		mem[  1687] = 11'd33;    
		mem[  1688] = 11'd23;    
		mem[  1689] = 11'd37;    
		mem[  1690] = 11'd27;    
		mem[  1691] = 11'd30;    
		mem[  1692] = 11'd66;    
		mem[  1693] = 11'd26;    
		mem[  1694] = 11'd65;    
		mem[  1695] = 11'd31;    
		mem[  1696] = 11'd60;    
		mem[  1697] = 11'd31;    
		mem[  1698] = 11'd22;    
		mem[  1699] = 11'd41;    
		mem[  1700] = 11'd24;    
		mem[  1701] = 11'd30;    
		mem[  1702] = 11'd32;    
		mem[  1703] = 11'd36;    
		mem[  1704] = 11'd25;    
		mem[  1705] = 11'd33;    
		mem[  1706] = 11'd32;    
		mem[  1707] = 11'd29;    
		mem[  1708] = 11'd26;    
		mem[  1709] = 11'd39;    
		mem[  1710] = 11'd28;    
		mem[  1711] = 11'd24;    
		mem[  1712] = 11'd40;    
		mem[  1713] = 11'd21;    
		mem[  1714] = 11'd33;    
		mem[  1715] = 11'd35;    
		mem[  1716] = 11'd33;    
		mem[  1717] = 11'd25;    
		mem[  1718] = 11'd36;    
		mem[  1719] = 11'd28;    
		mem[  1720] = 11'd29;    
		mem[  1721] = 11'd30;    
		mem[  1722] = 11'd37;    
		mem[  1723] = 11'd26;    
		mem[  1724] = 11'd29;    
		mem[  1725] = 11'd35;    
		mem[  1726] = 11'd31;    
		mem[  1727] = 11'd25;    
		mem[  1728] = 11'd33;    
		mem[  1729] = 11'd30;    
		mem[  1730] = 11'd24;    
		mem[  1731] = 11'd34;    
		mem[  1732] = 11'd27;    
		mem[  1733] = 11'd28;    
		mem[  1734] = 11'd27;    
		mem[  1735] = 11'd35;    
		mem[  1736] = 11'd27;    
		mem[  1737] = 11'd24;    
		mem[  1738] = 11'd36;    
		mem[  1739] = 11'd24;    
		mem[  1740] = 11'd29;    
		mem[  1741] = 11'd29;    
		mem[  1742] = 11'd33;    
		mem[  1743] = 11'd26;    
		mem[  1744] = 11'd27;    
		mem[  1745] = 11'd34;    
		mem[  1746] = 11'd26;    
		mem[  1747] = 11'd27;    
		mem[  1748] = 11'd31;    
		mem[  1749] = 11'd32;    
		mem[  1750] = 11'd25;    
		mem[  1751] = 11'd30;    
		mem[  1752] = 11'd31;    
		mem[  1753] = 11'd29;    
		mem[  1754] = 11'd25;    
		mem[  1755] = 11'd33;    
		mem[  1756] = 11'd29;    
		mem[  1757] = 11'd25;    
		mem[  1758] = 11'd33;    
		mem[  1759] = 11'd27;    
		mem[  1760] = 11'd29;    
		mem[  1761] = 11'd27;    
		mem[  1762] = 11'd34;    
		mem[  1763] = 11'd27;    
		mem[  1764] = 11'd25;    
		mem[  1765] = 11'd34;    
		mem[  1766] = 11'd26;    
		mem[  1767] = 11'd29;    
		mem[  1768] = 11'd29;    
		mem[  1769] = 11'd32;    
		mem[  1770] = 11'd27;    
		mem[  1771] = 11'd28;    
		mem[  1772] = 11'd32;    
		mem[  1773] = 11'd27;    
		mem[  1774] = 11'd28;    
		mem[  1775] = 11'd30;    
		mem[  1776] = 11'd31;    
		mem[  1777] = 11'd26;    
		mem[  1778] = 11'd28;    
		mem[  1779] = 11'd29;    
		mem[  1780] = 11'd26;    
		mem[  1781] = 11'd26;    
		mem[  1782] = 11'd28;    
		mem[  1783] = 11'd29;    
		mem[  1784] = 11'd26;    
		mem[  1785] = 11'd27;    
		mem[  1786] = 11'd29;    
		mem[  1787] = 11'd25;    
		mem[  1788] = 11'd27;    
		mem[  1789] = 11'd28;    
		mem[  1790] = 11'd30;    
		mem[  1791] = 11'd25;    
		mem[  1792] = 11'd26;    
		mem[  1793] = 11'd30;    
		mem[  1794] = 11'd25;    
		mem[  1795] = 11'd28;    
		mem[  1796] = 11'd27;    
		mem[  1797] = 11'd29;    
		mem[  1798] = 11'd27;    
		mem[  1799] = 11'd25;    
		mem[  1800] = 11'd30;    
		mem[  1801] = 11'd26;    
		mem[  1802] = 11'd27;    
		mem[  1803] = 11'd27;    
		mem[  1804] = 11'd29;    
		mem[  1805] = 11'd27;    
		mem[  1806] = 11'd26;    
		mem[  1807] = 11'd29;    
		mem[  1808] = 11'd27;    
		mem[  1809] = 11'd27;    
		mem[  1810] = 11'd26;    
		mem[  1811] = 11'd29;    
		mem[  1812] = 11'd28;    
		mem[  1813] = 11'd25;    
		mem[  1814] = 11'd29;    
		mem[  1815] = 11'd27;    
		mem[  1816] = 11'd28;    
		mem[  1817] = 11'd25;    
		mem[  1818] = 11'd29;    
		mem[  1819] = 11'd28;    
		mem[  1820] = 11'd26;    
		mem[  1821] = 11'd27;    
		mem[  1822] = 11'd28;    
		mem[  1823] = 11'd27;    
		mem[  1824] = 11'd27;    
		mem[  1825] = 11'd28;    
		mem[  1826] = 11'd28;    
		mem[  1827] = 11'd26;    
		mem[  1828] = 11'd27;    
		mem[  1829] = 11'd29;    
		mem[  1830] = 11'd26;    
		mem[  1831] = 11'd183;    
		mem[  1832] = 11'd30;    
		mem[  1833] = 11'd106;    
		mem[  1834] = 11'd68;    
		mem[  1835] = 11'd132;    
		mem[  1836] = 11'd192;    
		mem[  1837] = 11'd532;    
		mem[  1838] = 11'd244;    
		mem[  1839] = 11'd57;    
		mem[  1840] = 11'd24;    
		mem[  1841] = 11'd23;    
		mem[  1842] = 11'd35;    
		mem[  1843] = 11'd23;    
		mem[  1844] = 11'd58;    
		mem[  1845] = 11'd18;    
		mem[  1846] = 11'd28;    
		mem[  1847] = 11'd32;    
		mem[  1848] = 11'd30;    
		mem[  1849] = 11'd21;    
		mem[  1850] = 11'd32;    
		mem[  1851] = 11'd25;    
		mem[  1852] = 11'd27;    
		mem[  1853] = 11'd59;    
		mem[  1854] = 11'd24;    
		mem[  1855] = 11'd57;    
		mem[  1856] = 11'd28;    
		mem[  1857] = 11'd20;    
		mem[  1858] = 11'd33;    
		mem[  1859] = 11'd28;    
		mem[  1860] = 11'd20;    
		mem[  1861] = 11'd36;    
		mem[  1862] = 11'd22;    
		mem[  1863] = 11'd27;    
		mem[  1864] = 11'd28;    
		mem[  1865] = 11'd32;    
		mem[  1866] = 11'd22;    
		mem[  1867] = 11'd30;    
		mem[  1868] = 11'd28;    
		mem[  1869] = 11'd26;    
		mem[  1870] = 11'd23;    
		mem[  1871] = 11'd35;    
		mem[  1872] = 11'd25;    
		mem[  1873] = 11'd22;    
		mem[  1874] = 11'd34;    
		mem[  1875] = 11'd25;    
		mem[  1876] = 11'd24;    
		mem[  1877] = 11'd31;    
		mem[  1878] = 11'd29;    
		mem[  1879] = 11'd22;    
		mem[  1880] = 11'd33;    
		mem[  1881] = 11'd24;    
		mem[  1882] = 11'd27;    
		mem[  1883] = 11'd27;    
		mem[  1884] = 11'd32;    
		mem[  1885] = 11'd24;    
		mem[  1886] = 11'd26;    
		mem[  1887] = 11'd30;    
		mem[  1888] = 11'd26;    
		mem[  1889] = 11'd21;    
		mem[  1890] = 11'd30;    
		mem[  1891] = 11'd27;    
		mem[  1892] = 11'd21;    
		mem[  1893] = 11'd30;    
		mem[  1894] = 11'd24;    
		mem[  1895] = 11'd26;    
		mem[  1896] = 11'd23;    
		mem[  1897] = 11'd31;    
		mem[  1898] = 11'd24;    
		mem[  1899] = 11'd22;    
		mem[  1900] = 11'd32;    
		mem[  1901] = 11'd22;    
		mem[  1902] = 11'd25;    
		mem[  1903] = 11'd26;    
		mem[  1904] = 11'd30;    
		mem[  1905] = 11'd23;    
		mem[  1906] = 11'd23;    
		mem[  1907] = 11'd31;    
		mem[  1908] = 11'd20;    
		mem[  1909] = 11'd27;    
		mem[  1910] = 11'd27;    
		mem[  1911] = 11'd29;    
		mem[  1912] = 11'd23;    
		mem[  1913] = 11'd25;    
		mem[  1914] = 11'd29;    
		mem[  1915] = 11'd26;    
		mem[  1916] = 11'd22;    
		mem[  1917] = 11'd29;    
		mem[  1918] = 11'd26;    
		mem[  1919] = 11'd22;    
		mem[  1920] = 11'd29;    
		mem[  1921] = 11'd25;    
		mem[  1922] = 11'd26;    
		mem[  1923] = 11'd23;    
		mem[  1924] = 11'd30;    
		mem[  1925] = 11'd25;    
		mem[  1926] = 11'd22;    
		mem[  1927] = 11'd31;    
		mem[  1928] = 11'd23;    
		mem[  1929] = 11'd25;    
		mem[  1930] = 11'd26;    
		mem[  1931] = 11'd28;    
		mem[  1932] = 11'd25;    
		mem[  1933] = 11'd24;    
		mem[  1934] = 11'd29;    
		mem[  1935] = 11'd24;    
		mem[  1936] = 11'd25;    
		mem[  1937] = 11'd26;    
		mem[  1938] = 11'd28;    
		mem[  1939] = 11'd24;    
		mem[  1940] = 11'd26;    
		mem[  1941] = 11'd27;    
		mem[  1942] = 11'd26;    
		mem[  1943] = 11'd23;    
		mem[  1944] = 11'd27;    
		mem[  1945] = 11'd25;    
		mem[  1946] = 11'd22;    
		mem[  1947] = 11'd26;    
		mem[  1948] = 11'd25;    
		mem[  1949] = 11'd25;    
		mem[  1950] = 11'd22;    
		mem[  1951] = 11'd26;    
		mem[  1952] = 11'd26;    
		mem[  1953] = 11'd22;    
		mem[  1954] = 11'd24;    
		mem[  1955] = 11'd27;    
		mem[  1956] = 11'd23;    
		mem[  1957] = 11'd23;    
		mem[  1958] = 11'd26;    
		mem[  1959] = 11'd26;    
		mem[  1960] = 11'd23;    
		mem[  1961] = 11'd24;    
		mem[  1962] = 11'd26;    
		mem[  1963] = 11'd23;    
		mem[  1964] = 11'd24;    
		mem[  1965] = 11'd25;    
		mem[  1966] = 11'd26;    
		mem[  1967] = 11'd23;    
		mem[  1968] = 11'd24;    
		mem[  1969] = 11'd26;    
		mem[  1970] = 11'd22;    
		mem[  1971] = 11'd25;    
		mem[  1972] = 11'd25;    
		mem[  1973] = 11'd26;    
		mem[  1974] = 11'd24;    
		mem[  1975] = 11'd23;    
		mem[  1976] = 11'd26;    
		mem[  1977] = 11'd23;    
		mem[  1978] = 11'd25;    
		mem[  1979] = 11'd24;    
		mem[  1980] = 11'd26;    
		mem[  1981] = 11'd24;    
		mem[  1982] = 11'd23;    
		mem[  1983] = 11'd26;    
		mem[  1984] = 11'd24;    
		mem[  1985] = 11'd24;    
		mem[  1986] = 11'd24;    
		mem[  1987] = 11'd26;    
		mem[  1988] = 11'd24;    
		mem[  1989] = 11'd24;    
		mem[  1990] = 11'd25;    
		mem[  1991] = 11'd25;    
		mem[  1992] = 11'd24;    
		mem[  1993] = 11'd24;    
		mem[  1994] = 11'd25;    
		mem[  1995] = 11'd25;    
		mem[  1996] = 11'd23;    
		mem[  1997] = 11'd25;    
		mem[  1998] = 11'd25;    
		mem[  1999] = 11'd25;    
		mem[  2000] = 11'd23;    
		mem[  2001] = 11'd25;    
		mem[  2002] = 11'd25;    
		mem[  2003] = 11'd193;    
		mem[  2004] = 11'd55;    
		mem[  2005] = 11'd1250;    
		mem[  2006] = 11'd44;    
		mem[  2007] = 11'd22;    
		mem[  2008] = 11'd17;    
		mem[  2009] = 11'd45;    
		mem[  2010] = 11'd16;    
		mem[  2011] = 11'd21;    
		mem[  2012] = 11'd44;    
		mem[  2013] = 11'd22;    
		mem[  2014] = 11'd16;    
		mem[  2015] = 11'd20;    
		mem[  2016] = 11'd26;    
		mem[  2017] = 11'd15;    
		mem[  2018] = 11'd21;    
		mem[  2019] = 11'd19;    
		mem[  2020] = 11'd25;    
		mem[  2021] = 11'd22;    
		mem[  2022] = 11'd16;    
		mem[  2023] = 11'd20;    
		mem[  2024] = 11'd26;    
		mem[  2025] = 11'd15;    
		mem[  2026] = 11'd21;    
		mem[  2027] = 11'd19;    
		mem[  2028] = 11'd25;    
		mem[  2029] = 11'd21;    
		mem[  2030] = 11'd17;    
		mem[  2031] = 11'd20;    
		mem[  2032] = 11'd25;    
		mem[  2033] = 11'd16;    
		mem[  2034] = 11'd21;    
		mem[  2035] = 11'd18;    
		mem[  2036] = 11'd26;    
		mem[  2037] = 11'd21;    
		mem[  2038] = 11'd17;    
		mem[  2039] = 11'd19;    
		mem[  2040] = 11'd26;    
		mem[  2041] = 11'd16;    
		mem[  2042] = 11'd21;    
		mem[  2043] = 11'd18;    
		mem[  2044] = 11'd25;    
		mem[  2045] = 11'd22;    
		mem[  2046] = 11'd16;    
		mem[  2047] = 11'd20;    
		mem[  2048] = 11'd25;    
		mem[  2049] = 11'd16;    
		mem[  2050] = 11'd21;    
		mem[  2051] = 11'd19;    
		mem[  2052] = 11'd25;    
		mem[  2053] = 11'd21;    
		mem[  2054] = 11'd17;    
		mem[  2055] = 11'd20;    
		mem[  2056] = 11'd25;    
		mem[  2057] = 11'd16;    
		mem[  2058] = 11'd21;    
		mem[  2059] = 11'd19;    
		mem[  2060] = 11'd25;    
		mem[  2061] = 11'd21;    
		mem[  2062] = 11'd17;    
		mem[  2063] = 11'd20;    
		mem[  2064] = 11'd25;    
		mem[  2065] = 11'd16;    
		mem[  2066] = 11'd21;    
		mem[  2067] = 11'd19;    
		mem[  2068] = 11'd24;    
		mem[  2069] = 11'd22;    
		mem[  2070] = 11'd17;    
		mem[  2071] = 11'd20;    
		mem[  2072] = 11'd24;    
		mem[  2073] = 11'd17;    
		mem[  2074] = 11'd21;    
		mem[  2075] = 11'd19;    
		mem[  2076] = 11'd24;    
		mem[  2077] = 11'd21;    
		mem[  2078] = 11'd18;    
		mem[  2079] = 11'd20;    
		mem[  2080] = 11'd24;    
		mem[  2081] = 11'd17;    
		mem[  2082] = 11'd21;    
		mem[  2083] = 11'd19;    
		mem[  2084] = 11'd24;    
		mem[  2085] = 11'd21;    
		mem[  2086] = 11'd18;    
		mem[  2087] = 11'd20;    
		mem[  2088] = 11'd24;    
		mem[  2089] = 11'd17;    
		mem[  2090] = 11'd21;    
		mem[  2091] = 11'd19;    
		mem[  2092] = 11'd24;    
		mem[  2093] = 11'd21;    
		mem[  2094] = 11'd17;    
		mem[  2095] = 11'd21;    
		mem[  2096] = 11'd24;    
		mem[  2097] = 11'd17;    
		mem[  2098] = 11'd21;    
		mem[  2099] = 11'd19;    
		mem[  2100] = 11'd23;    
		mem[  2101] = 11'd22;    
		mem[  2102] = 11'd17;    
		mem[  2103] = 11'd20;    
		mem[  2104] = 11'd24;    
		mem[  2105] = 11'd17;    
		mem[  2106] = 11'd21;    
		mem[  2107] = 11'd20;    
		mem[  2108] = 11'd23;    
		mem[  2109] = 11'd21;    
		mem[  2110] = 11'd18;    
		mem[  2111] = 11'd21;    
		mem[  2112] = 11'd23;    
		mem[  2113] = 11'd17;    
		mem[  2114] = 11'd21;    
		mem[  2115] = 11'd20;    
		mem[  2116] = 11'd23;    
		mem[  2117] = 11'd21;    
		mem[  2118] = 11'd18;    
		mem[  2119] = 11'd20;    
		mem[  2120] = 11'd24;    
		mem[  2121] = 11'd17;    
		mem[  2122] = 11'd21;    
		mem[  2123] = 11'd20;    
		mem[  2124] = 11'd23;    
		mem[  2125] = 11'd21;    
		mem[  2126] = 11'd18;    
		mem[  2127] = 11'd20;    
		mem[  2128] = 11'd23;    
		mem[  2129] = 11'd18;    
		mem[  2130] = 11'd21;    
		mem[  2131] = 11'd20;    
		mem[  2132] = 11'd23;    
		mem[  2133] = 11'd20;    
		mem[  2134] = 11'd19;    
		mem[  2135] = 11'd20;    
		mem[  2136] = 11'd23;    
		mem[  2137] = 11'd18;    
		mem[  2138] = 11'd21;    
		mem[  2139] = 11'd20;    
		mem[  2140] = 11'd22;    
		mem[  2141] = 11'd21;    
		mem[  2142] = 11'd19;    
		mem[  2143] = 11'd20;    
		mem[  2144] = 11'd55;    
		mem[  2145] = 11'd83;    
		mem[  2146] = 11'd65;    
		mem[  2147] = 11'd20;    
		mem[  2148] = 11'd83;    
		mem[  2149] = 11'd61;    
		mem[  2150] = 11'd22;    
		mem[  2151] = 11'd80;    
		mem[  2152] = 11'd62;    
		mem[  2153] = 11'd21;    
		mem[  2154] = 11'd81;    
		mem[  2155] = 11'd62;    
		mem[  2156] = 11'd22;    
		mem[  2157] = 11'd78;    
		mem[  2158] = 11'd63;    
		mem[  2159] = 11'd21;    
		mem[  2160] = 11'd82;    
		mem[  2161] = 11'd61;    
		mem[  2162] = 11'd21;    
		mem[  2163] = 11'd79;    
		mem[  2164] = 11'd63;    
		mem[  2165] = 11'd21;    
		mem[  2166] = 11'd83;    
		mem[  2167] = 11'd60;    
		mem[  2168] = 11'd22;    
		mem[  2169] = 11'd80;    
		mem[  2170] = 11'd60;    
		mem[  2171] = 11'd20;    
		mem[  2172] = 11'd86;    
		mem[  2173] = 11'd61;    
		mem[  2174] = 11'd21;    
		mem[  2175] = 11'd80;    
		mem[  2176] = 11'd58;    
		mem[  2177] = 11'd108;    
		mem[  2178] = 11'd62;    
		mem[  2179] = 11'd20;    
		mem[  2180] = 11'd78;    
		mem[  2181] = 11'd64;    
		mem[  2182] = 11'd19;    

	end
	
endmodule

