module pacman_intermission_converted(in, out, clk); //ok
	 input [11:0] in;
	 input clk;
	 output reg [8:0] out;
	 
	 reg  [8:0] mem [0:2838];
	 always @(posedge clk) out  =  mem[ in ];
	 
	 initial begin
		mem[     0] = 9'd91;    
		mem[     1] = 9'd31;    
		mem[     2] = 9'd61;    
		mem[     3] = 9'd22;    
		mem[     4] = 9'd113;    
		mem[     5] = 9'd65;    
		mem[     6] = 9'd33;    
		mem[     7] = 9'd33;    
		mem[     8] = 9'd63;    
		mem[     9] = 9'd64;    
		mem[    10] = 9'd68;    
		mem[    11] = 9'd28;    
		mem[    12] = 9'd33;    
		mem[    13] = 9'd68;    
		mem[    14] = 9'd32;    
		mem[    15] = 9'd25;    
		mem[    16] = 9'd65;    
		mem[    17] = 9'd58;    
		mem[    18] = 9'd65;    
		mem[    19] = 9'd58;    
		mem[    20] = 9'd64;    
		mem[    21] = 9'd59;    
		mem[    22] = 9'd64;    
		mem[    23] = 9'd58;    
		mem[    24] = 9'd64;    
		mem[    25] = 9'd59;    
		mem[    26] = 9'd64;    
		mem[    27] = 9'd32;    
		mem[    28] = 9'd26;    
		mem[    29] = 9'd64;    
		mem[    30] = 9'd59;    
		mem[    31] = 9'd64;    
		mem[    32] = 9'd32;    
		mem[    33] = 9'd26;    
		mem[    34] = 9'd64;    
		mem[    35] = 9'd59;    
		mem[    36] = 9'd64;    
		mem[    37] = 9'd32;    
		mem[    38] = 9'd26;    
		mem[    39] = 9'd31;    
		mem[    40] = 9'd33;    
		mem[    41] = 9'd59;    
		mem[    42] = 9'd64;    
		mem[    43] = 9'd32;    
		mem[    44] = 9'd27;    
		mem[    45] = 9'd30;    
		mem[    46] = 9'd33;    
		mem[    47] = 9'd60;    
		mem[    48] = 9'd63;    
		mem[    49] = 9'd32;    
		mem[    50] = 9'd27;    
		mem[    51] = 9'd31;    
		mem[    52] = 9'd32;    
		mem[    53] = 9'd60;    
		mem[    54] = 9'd63;    
		mem[    55] = 9'd32;    
		mem[    56] = 9'd27;    
		mem[    57] = 9'd31;    
		mem[    58] = 9'd32;    
		mem[    59] = 9'd60;    
		mem[    60] = 9'd60;    
		mem[    61] = 9'd62;    
		mem[    62] = 9'd31;    
		mem[    63] = 9'd31;    
		mem[    64] = 9'd32;    
		mem[    65] = 9'd30;    
		mem[    66] = 9'd31;    
		mem[    67] = 9'd30;    
		mem[    68] = 9'd31;    
		mem[    69] = 9'd30;    
		mem[    70] = 9'd32;    
		mem[    71] = 9'd30;    
		mem[    72] = 9'd31;    
		mem[    73] = 9'd30;    
		mem[    74] = 9'd31;    
		mem[    75] = 9'd30;    
		mem[    76] = 9'd32;    
		mem[    77] = 9'd29;    
		mem[    78] = 9'd32;    
		mem[    79] = 9'd29;    
		mem[    80] = 9'd32;    
		mem[    81] = 9'd30;    
		mem[    82] = 9'd32;    
		mem[    83] = 9'd32;    
		mem[    84] = 9'd33;    
		mem[    85] = 9'd31;    
		mem[    86] = 9'd34;    
		mem[    87] = 9'd32;    
		mem[    88] = 9'd33;    
		mem[    89] = 9'd31;    
		mem[    90] = 9'd34;    
		mem[    91] = 9'd31;    
		mem[    92] = 9'd34;    
		mem[    93] = 9'd32;    
		mem[    94] = 9'd33;    
		mem[    95] = 9'd31;    
		mem[    96] = 9'd33;    
		mem[    97] = 9'd32;    
		mem[    98] = 9'd34;    
		mem[    99] = 9'd31;    
		mem[   100] = 9'd34;    
		mem[   101] = 9'd31;    
		mem[   102] = 9'd33;    
		mem[   103] = 9'd32;    
		mem[   104] = 9'd33;    
		mem[   105] = 9'd30;    
		mem[   106] = 9'd31;    
		mem[   107] = 9'd30;    
		mem[   108] = 9'd31;    
		mem[   109] = 9'd31;    
		mem[   110] = 9'd31;    
		mem[   111] = 9'd30;    
		mem[   112] = 9'd31;    
		mem[   113] = 9'd30;    
		mem[   114] = 9'd31;    
		mem[   115] = 9'd31;    
		mem[   116] = 9'd31;    
		mem[   117] = 9'd30;    
		mem[   118] = 9'd31;    
		mem[   119] = 9'd30;    
		mem[   120] = 9'd31;    
		mem[   121] = 9'd30;    
		mem[   122] = 9'd32;    
		mem[   123] = 9'd30;    
		mem[   124] = 9'd31;    
		mem[   125] = 9'd30;    
		mem[   126] = 9'd31;    
		mem[   127] = 9'd30;    
		mem[   128] = 9'd33;    
		mem[   129] = 9'd88;    
		mem[   130] = 9'd65;    
		mem[   131] = 9'd58;    
		mem[   132] = 9'd64;    
		mem[   133] = 9'd32;    
		mem[   134] = 9'd25;    
		mem[   135] = 9'd66;    
		mem[   136] = 9'd58;    
		mem[   137] = 9'd64;    
		mem[   138] = 9'd58;    
		mem[   139] = 9'd65;    
		mem[   140] = 9'd58;    
		mem[   141] = 9'd64;    
		mem[   142] = 9'd58;    
		mem[   143] = 9'd65;    
		mem[   144] = 9'd58;    
		mem[   145] = 9'd65;    
		mem[   146] = 9'd57;    
		mem[   147] = 9'd65;    
		mem[   148] = 9'd58;    
		mem[   149] = 9'd64;    
		mem[   150] = 9'd59;    
		mem[   151] = 9'd64;    
		mem[   152] = 9'd59;    
		mem[   153] = 9'd61;    
		mem[   154] = 9'd30;    
		mem[   155] = 9'd32;    
		mem[   156] = 9'd30;    
		mem[   157] = 9'd31;    
		mem[   158] = 9'd32;    
		mem[   159] = 9'd30;    
		mem[   160] = 9'd31;    
		mem[   161] = 9'd30;    
		mem[   162] = 9'd32;    
		mem[   163] = 9'd30;    
		mem[   164] = 9'd31;    
		mem[   165] = 9'd30;    
		mem[   166] = 9'd31;    
		mem[   167] = 9'd30;    
		mem[   168] = 9'd31;    
		mem[   169] = 9'd30;    
		mem[   170] = 9'd32;    
		mem[   171] = 9'd30;    
		mem[   172] = 9'd31;    
		mem[   173] = 9'd30;    
		mem[   174] = 9'd31;    
		mem[   175] = 9'd30;    
		mem[   176] = 9'd36;    
		mem[   177] = 9'd64;    
		mem[   178] = 9'd15;    
		mem[   179] = 9'd79;    
		mem[   180] = 9'd33;    
		mem[   181] = 9'd99;    
		mem[   182] = 9'd28;    
		mem[   183] = 9'd34;    
		mem[   184] = 9'd58;    
		mem[   185] = 9'd22;    
		mem[   186] = 9'd50;    
		mem[   187] = 9'd67;    
		mem[   188] = 9'd66;    
		mem[   189] = 9'd32;    
		mem[   190] = 9'd32;    
		mem[   191] = 9'd62;    
		mem[   192] = 9'd61;    
		mem[   193] = 9'd63;    
		mem[   194] = 9'd29;    
		mem[   195] = 9'd30;    
		mem[   196] = 9'd62;    
		mem[   197] = 9'd61;    
		mem[   198] = 9'd63;    
		mem[   199] = 9'd29;    
		mem[   200] = 9'd30;    
		mem[   201] = 9'd62;    
		mem[   202] = 9'd61;    
		mem[   203] = 9'd63;    
		mem[   204] = 9'd29;    
		mem[   205] = 9'd31;    
		mem[   206] = 9'd61;    
		mem[   207] = 9'd61;    
		mem[   208] = 9'd63;    
		mem[   209] = 9'd14;    
		mem[   210] = 9'd15;    
		mem[   211] = 9'd31;    
		mem[   212] = 9'd61;    
		mem[   213] = 9'd61;    
		mem[   214] = 9'd63;    
		mem[   215] = 9'd14;    
		mem[   216] = 9'd15;    
		mem[   217] = 9'd31;    
		mem[   218] = 9'd61;    
		mem[   219] = 9'd61;    
		mem[   220] = 9'd63;    
		mem[   221] = 9'd14;    
		mem[   222] = 9'd15;    
		mem[   223] = 9'd31;    
		mem[   224] = 9'd61;    
		mem[   225] = 9'd61;    
		mem[   226] = 9'd63;    
		mem[   227] = 9'd29;    
		mem[   228] = 9'd31;    
		mem[   229] = 9'd62;    
		mem[   230] = 9'd60;    
		mem[   231] = 9'd63;    
		mem[   232] = 9'd30;    
		mem[   233] = 9'd30;    
		mem[   234] = 9'd62;    
		mem[   235] = 9'd61;    
		mem[   236] = 9'd62;    
		mem[   237] = 9'd30;    
		mem[   238] = 9'd33;    
		mem[   239] = 9'd59;    
		mem[   240] = 9'd32;    
		mem[   241] = 9'd29;    
		mem[   242] = 9'd31;    
		mem[   243] = 9'd30;    
		mem[   244] = 9'd31;    
		mem[   245] = 9'd30;    
		mem[   246] = 9'd30;    
		mem[   247] = 9'd31;    
		mem[   248] = 9'd30;    
		mem[   249] = 9'd31;    
		mem[   250] = 9'd30;    
		mem[   251] = 9'd31;    
		mem[   252] = 9'd31;    
		mem[   253] = 9'd31;    
		mem[   254] = 9'd30;    
		mem[   255] = 9'd31;    
		mem[   256] = 9'd31;    
		mem[   257] = 9'd30;    
		mem[   258] = 9'd31;    
		mem[   259] = 9'd31;    
		mem[   260] = 9'd31;    
		mem[   261] = 9'd32;    
		mem[   262] = 9'd40;    
		mem[   263] = 9'd38;    
		mem[   264] = 9'd40;    
		mem[   265] = 9'd38;    
		mem[   266] = 9'd39;    
		mem[   267] = 9'd39;    
		mem[   268] = 9'd39;    
		mem[   269] = 9'd39;    
		mem[   270] = 9'd39;    
		mem[   271] = 9'd38;    
		mem[   272] = 9'd40;    
		mem[   273] = 9'd38;    
		mem[   274] = 9'd39;    
		mem[   275] = 9'd39;    
		mem[   276] = 9'd39;    
		mem[   277] = 9'd38;    
		mem[   278] = 9'd40;    
		mem[   279] = 9'd38;    
		mem[   280] = 9'd40;    
		mem[   281] = 9'd35;    
		mem[   282] = 9'd37;    
		mem[   283] = 9'd35;    
		mem[   284] = 9'd37;    
		mem[   285] = 9'd36;    
		mem[   286] = 9'd38;    
		mem[   287] = 9'd36;    
		mem[   288] = 9'd37;    
		mem[   289] = 9'd36;    
		mem[   290] = 9'd37;    
		mem[   291] = 9'd36;    
		mem[   292] = 9'd37;    
		mem[   293] = 9'd36;    
		mem[   294] = 9'd37;    
		mem[   295] = 9'd36;    
		mem[   296] = 9'd38;    
		mem[   297] = 9'd36;    
		mem[   298] = 9'd37;    
		mem[   299] = 9'd36;    
		mem[   300] = 9'd144;    
		mem[   301] = 9'd77;    
		mem[   302] = 9'd39;    
		mem[   303] = 9'd15;    
		mem[   304] = 9'd15;    
		mem[   305] = 9'd78;    
		mem[   306] = 9'd73;    
		mem[   307] = 9'd35;    
		mem[   308] = 9'd36;    
		mem[   309] = 9'd76;    
		mem[   310] = 9'd37;    
		mem[   311] = 9'd16;    
		mem[   312] = 9'd87;    
		mem[   313] = 9'd21;    
		mem[   314] = 9'd64;    
		mem[   315] = 9'd78;    
		mem[   316] = 9'd82;    
		mem[   317] = 9'd21;    
		mem[   318] = 9'd65;    
		mem[   319] = 9'd78;    
		mem[   320] = 9'd81;    
		mem[   321] = 9'd21;    
		mem[   322] = 9'd65;    
		mem[   323] = 9'd46;    
		mem[   324] = 9'd21;    
		mem[   325] = 9'd12;    
		mem[   326] = 9'd81;    
		mem[   327] = 9'd84;    
		mem[   328] = 9'd41;    
		mem[   329] = 9'd42;    
		mem[   330] = 9'd42;    
		mem[   331] = 9'd40;    
		mem[   332] = 9'd43;    
		mem[   333] = 9'd39;    
		mem[   334] = 9'd43;    
		mem[   335] = 9'd39;    
		mem[   336] = 9'd43;    
		mem[   337] = 9'd39;    
		mem[   338] = 9'd42;    
		mem[   339] = 9'd40;    
		mem[   340] = 9'd42;    
		mem[   341] = 9'd40;    
		mem[   342] = 9'd42;    
		mem[   343] = 9'd57;    
		mem[   344] = 9'd12;    
		mem[   345] = 9'd30;    
		mem[   346] = 9'd63;    
		mem[   347] = 9'd60;    
		mem[   348] = 9'd34;    
		mem[   349] = 9'd14;    
		mem[   350] = 9'd13;    
		mem[   351] = 9'd60;    
		mem[   352] = 9'd64;    
		mem[   353] = 9'd60;    
		mem[   354] = 9'd34;    
		mem[   355] = 9'd14;    
		mem[   356] = 9'd13;    
		mem[   357] = 9'd60;    
		mem[   358] = 9'd64;    
		mem[   359] = 9'd60;    
		mem[   360] = 9'd34;    
		mem[   361] = 9'd14;    
		mem[   362] = 9'd13;    
		mem[   363] = 9'd60;    
		mem[   364] = 9'd64;    
		mem[   365] = 9'd60;    
		mem[   366] = 9'd34;    
		mem[   367] = 9'd14;    
		mem[   368] = 9'd13;    
		mem[   369] = 9'd60;    
		mem[   370] = 9'd64;    
		mem[   371] = 9'd60;    
		mem[   372] = 9'd34;    
		mem[   373] = 9'd14;    
		mem[   374] = 9'd13;    
		mem[   375] = 9'd60;    
		mem[   376] = 9'd63;    
		mem[   377] = 9'd61;    
		mem[   378] = 9'd34;    
		mem[   379] = 9'd14;    
		mem[   380] = 9'd32;    
		mem[   381] = 9'd115;    
		mem[   382] = 9'd91;    
		mem[   383] = 9'd32;    
		mem[   384] = 9'd121;    
		mem[   385] = 9'd92;    
		mem[   386] = 9'd32;    
		mem[   387] = 9'd121;    
		mem[   388] = 9'd93;    
		mem[   389] = 9'd7;    
		mem[   390] = 9'd65;    
		mem[   391] = 9'd35;    
		mem[   392] = 9'd29;    
		mem[   393] = 9'd60;    
		mem[   394] = 9'd60;    
		mem[   395] = 9'd31;    
		mem[   396] = 9'd31;    
		mem[   397] = 9'd63;    
		mem[   398] = 9'd28;    
		mem[   399] = 9'd32;    
		mem[   400] = 9'd35;    
		mem[   401] = 9'd25;    
		mem[   402] = 9'd32;    
		mem[   403] = 9'd18;    
		mem[   404] = 9'd12;    
		mem[   405] = 9'd35;    
		mem[   406] = 9'd28;    
		mem[   407] = 9'd29;    
		mem[   408] = 9'd31;    
		mem[   409] = 9'd34;    
		mem[   410] = 9'd30;    
		mem[   411] = 9'd60;    
		mem[   412] = 9'd31;    
		mem[   413] = 9'd30;    
		mem[   414] = 9'd31;    
		mem[   415] = 9'd29;    
		mem[   416] = 9'd31;    
		mem[   417] = 9'd31;    
		mem[   418] = 9'd30;    
		mem[   419] = 9'd31;    
		mem[   420] = 9'd30;    
		mem[   421] = 9'd31;    
		mem[   422] = 9'd30;    
		mem[   423] = 9'd31;    
		mem[   424] = 9'd31;    
		mem[   425] = 9'd31;    
		mem[   426] = 9'd30;    
		mem[   427] = 9'd31;    
		mem[   428] = 9'd31;    
		mem[   429] = 9'd30;    
		mem[   430] = 9'd31;    
		mem[   431] = 9'd31;    
		mem[   432] = 9'd30;    
		mem[   433] = 9'd31;    
		mem[   434] = 9'd31;    
		mem[   435] = 9'd30;    
		mem[   436] = 9'd31;    
		mem[   437] = 9'd31;    
		mem[   438] = 9'd31;    
		mem[   439] = 9'd30;    
		mem[   440] = 9'd31;    
		mem[   441] = 9'd30;    
		mem[   442] = 9'd31;    
		mem[   443] = 9'd30;    
		mem[   444] = 9'd31;    
		mem[   445] = 9'd30;    
		mem[   446] = 9'd32;    
		mem[   447] = 9'd30;    
		mem[   448] = 9'd31;    
		mem[   449] = 9'd30;    
		mem[   450] = 9'd31;    
		mem[   451] = 9'd30;    
		mem[   452] = 9'd32;    
		mem[   453] = 9'd30;    
		mem[   454] = 9'd31;    
		mem[   455] = 9'd30;    
		mem[   456] = 9'd32;    
		mem[   457] = 9'd30;    
		mem[   458] = 9'd31;    
		mem[   459] = 9'd30;    
		mem[   460] = 9'd31;    
		mem[   461] = 9'd30;    
		mem[   462] = 9'd31;    
		mem[   463] = 9'd30;    
		mem[   464] = 9'd31;    
		mem[   465] = 9'd30;    
		mem[   466] = 9'd31;    
		mem[   467] = 9'd31;    
		mem[   468] = 9'd30;    
		mem[   469] = 9'd31;    
		mem[   470] = 9'd31;    
		mem[   471] = 9'd30;    
		mem[   472] = 9'd31;    
		mem[   473] = 9'd30;    
		mem[   474] = 9'd31;    
		mem[   475] = 9'd31;    
		mem[   476] = 9'd30;    
		mem[   477] = 9'd31;    
		mem[   478] = 9'd31;    
		mem[   479] = 9'd30;    
		mem[   480] = 9'd27;    
		mem[   481] = 9'd28;    
		mem[   482] = 9'd105;    
		mem[   483] = 9'd23;    
		mem[   484] = 9'd80;    
		mem[   485] = 9'd49;    
		mem[   486] = 9'd52;    
		mem[   487] = 9'd53;    
		mem[   488] = 9'd50;    
		mem[   489] = 9'd52;    
		mem[   490] = 9'd30;    
		mem[   491] = 9'd20;    
		mem[   492] = 9'd55;    
		mem[   493] = 9'd50;    
		mem[   494] = 9'd53;    
		mem[   495] = 9'd46;    
		mem[   496] = 9'd27;    
		mem[   497] = 9'd23;    
		mem[   498] = 9'd52;    
		mem[   499] = 9'd47;    
		mem[   500] = 9'd51;    
		mem[   501] = 9'd44;    
		mem[   502] = 9'd28;    
		mem[   503] = 9'd22;    
		mem[   504] = 9'd53;    
		mem[   505] = 9'd47;    
		mem[   506] = 9'd50;    
		mem[   507] = 9'd46;    
		mem[   508] = 9'd26;    
		mem[   509] = 9'd23;    
		mem[   510] = 9'd52;    
		mem[   511] = 9'd47;    
		mem[   512] = 9'd51;    
		mem[   513] = 9'd49;    
		mem[   514] = 9'd26;    
		mem[   515] = 9'd22;    
		mem[   516] = 9'd25;    
		mem[   517] = 9'd24;    
		mem[   518] = 9'd25;    
		mem[   519] = 9'd23;    
		mem[   520] = 9'd25;    
		mem[   521] = 9'd24;    
		mem[   522] = 9'd25;    
		mem[   523] = 9'd24;    
		mem[   524] = 9'd24;    
		mem[   525] = 9'd25;    
		mem[   526] = 9'd24;    
		mem[   527] = 9'd25;    
		mem[   528] = 9'd24;    
		mem[   529] = 9'd25;    
		mem[   530] = 9'd24;    
		mem[   531] = 9'd25;    
		mem[   532] = 9'd24;    
		mem[   533] = 9'd25;    
		mem[   534] = 9'd24;    
		mem[   535] = 9'd25;    
		mem[   536] = 9'd24;    
		mem[   537] = 9'd25;    
		mem[   538] = 9'd24;    
		mem[   539] = 9'd25;    
		mem[   540] = 9'd24;    
		mem[   541] = 9'd25;    
		mem[   542] = 9'd23;    
		mem[   543] = 9'd26;    
		mem[   544] = 9'd98;    
		mem[   545] = 9'd50;    
		mem[   546] = 9'd25;    
		mem[   547] = 9'd24;    
		mem[   548] = 9'd47;    
		mem[   549] = 9'd50;    
		mem[   550] = 9'd50;    
		mem[   551] = 9'd25;    
		mem[   552] = 9'd24;    
		mem[   553] = 9'd47;    
		mem[   554] = 9'd50;    
		mem[   555] = 9'd50;    
		mem[   556] = 9'd24;    
		mem[   557] = 9'd25;    
		mem[   558] = 9'd46;    
		mem[   559] = 9'd50;    
		mem[   560] = 9'd50;    
		mem[   561] = 9'd25;    
		mem[   562] = 9'd24;    
		mem[   563] = 9'd47;    
		mem[   564] = 9'd50;    
		mem[   565] = 9'd50;    
		mem[   566] = 9'd25;    
		mem[   567] = 9'd24;    
		mem[   568] = 9'd47;    
		mem[   569] = 9'd50;    
		mem[   570] = 9'd49;    
		mem[   571] = 9'd25;    
		mem[   572] = 9'd25;    
		mem[   573] = 9'd47;    
		mem[   574] = 9'd50;    
		mem[   575] = 9'd49;    
		mem[   576] = 9'd25;    
		mem[   577] = 9'd24;    
		mem[   578] = 9'd47;    
		mem[   579] = 9'd49;    
		mem[   580] = 9'd24;    
		mem[   581] = 9'd25;    
		mem[   582] = 9'd25;    
		mem[   583] = 9'd24;    
		mem[   584] = 9'd25;    
		mem[   585] = 9'd24;    
		mem[   586] = 9'd26;    
		mem[   587] = 9'd24;    
		mem[   588] = 9'd24;    
		mem[   589] = 9'd24;    
		mem[   590] = 9'd26;    
		mem[   591] = 9'd23;    
		mem[   592] = 9'd75;    
		mem[   593] = 9'd22;    
		mem[   594] = 9'd49;    
		mem[   595] = 9'd24;    
		mem[   596] = 9'd76;    
		mem[   597] = 9'd48;    
		mem[   598] = 9'd27;    
		mem[   599] = 9'd10;    
		mem[   600] = 9'd14;    
		mem[   601] = 9'd46;    
		mem[   602] = 9'd50;    
		mem[   603] = 9'd50;    
		mem[   604] = 9'd23;    
		mem[   605] = 9'd24;    
		mem[   606] = 9'd51;    
		mem[   607] = 9'd46;    
		mem[   608] = 9'd52;    
		mem[   609] = 9'd37;    
		mem[   610] = 9'd8;    
		mem[   611] = 9'd53;    
		mem[   612] = 9'd24;    
		mem[   613] = 9'd72;    
		mem[   614] = 9'd25;    
		mem[   615] = 9'd75;    
		mem[   616] = 9'd20;    
		mem[   617] = 9'd26;    
		mem[   618] = 9'd46;    
		mem[   619] = 9'd14;    
		mem[   620] = 9'd38;    
		mem[   621] = 9'd50;    
		mem[   622] = 9'd50;    
		mem[   623] = 9'd24;    
		mem[   624] = 9'd24;    
		mem[   625] = 9'd49;    
		mem[   626] = 9'd48;    
		mem[   627] = 9'd51;    
		mem[   628] = 9'd47;    
		mem[   629] = 9'd48;    
		mem[   630] = 9'd50;    
		mem[   631] = 9'd24;    
		mem[   632] = 9'd25;    
		mem[   633] = 9'd25;    
		mem[   634] = 9'd24;    
		mem[   635] = 9'd25;    
		mem[   636] = 9'd24;    
		mem[   637] = 9'd25;    
		mem[   638] = 9'd24;    
		mem[   639] = 9'd25;    
		mem[   640] = 9'd24;    
		mem[   641] = 9'd25;    
		mem[   642] = 9'd25;    
		mem[   643] = 9'd49;    
		mem[   644] = 9'd71;    
		mem[   645] = 9'd25;    
		mem[   646] = 9'd52;    
		mem[   647] = 9'd24;    
		mem[   648] = 9'd71;    
		mem[   649] = 9'd24;    
		mem[   650] = 9'd75;    
		mem[   651] = 9'd50;    
		mem[   652] = 9'd23;    
		mem[   653] = 9'd24;    
		mem[   654] = 9'd50;    
		mem[   655] = 9'd46;    
		mem[   656] = 9'd52;    
		mem[   657] = 9'd24;    
		mem[   658] = 9'd87;    
		mem[   659] = 9'd65;    
		mem[   660] = 9'd23;    
		mem[   661] = 9'd86;    
		mem[   662] = 9'd65;    
		mem[   663] = 9'd23;    
		mem[   664] = 9'd86;    
		mem[   665] = 9'd66;    
		mem[   666] = 9'd22;    
		mem[   667] = 9'd87;    
		mem[   668] = 9'd65;    
		mem[   669] = 9'd22;    
		mem[   670] = 9'd247;    
		mem[   671] = 9'd264;    
		mem[   672] = 9'd21;    
		mem[   673] = 9'd82;    
		mem[   674] = 9'd62;    
		mem[   675] = 9'd21;    
		mem[   676] = 9'd82;    
		mem[   677] = 9'd63;    
		mem[   678] = 9'd21;    
		mem[   679] = 9'd80;    
		mem[   680] = 9'd63;    
		mem[   681] = 9'd21;    
		mem[   682] = 9'd79;    
		mem[   683] = 9'd63;    
		mem[   684] = 9'd22;    
		mem[   685] = 9'd79;    
		mem[   686] = 9'd63;    
		mem[   687] = 9'd20;    
		mem[   688] = 9'd81;    
		mem[   689] = 9'd61;    
		mem[   690] = 9'd22;    
		mem[   691] = 9'd81;    
		mem[   692] = 9'd61;    
		mem[   693] = 9'd21;    
		mem[   694] = 9'd82;    
		mem[   695] = 9'd61;    
		mem[   696] = 9'd21;    
		mem[   697] = 9'd245;    
		mem[   698] = 9'd208;    
		mem[   699] = 9'd67;    
		mem[   700] = 9'd30;    
		mem[   701] = 9'd33;    
		mem[   702] = 9'd68;    
		mem[   703] = 9'd61;    
		mem[   704] = 9'd69;    
		mem[   705] = 9'd61;    
		mem[   706] = 9'd70;    
		mem[   707] = 9'd32;    
		mem[   708] = 9'd15;    
		mem[   709] = 9'd80;    
		mem[   710] = 9'd33;    
		mem[   711] = 9'd98;    
		mem[   712] = 9'd28;    
		mem[   713] = 9'd29;    
		mem[   714] = 9'd63;    
		mem[   715] = 9'd31;    
		mem[   716] = 9'd94;    
		mem[   717] = 9'd28;    
		mem[   718] = 9'd29;    
		mem[   719] = 9'd63;    
		mem[   720] = 9'd31;    
		mem[   721] = 9'd28;    
		mem[   722] = 9'd66;    
		mem[   723] = 9'd28;    
		mem[   724] = 9'd29;    
		mem[   725] = 9'd63;    
		mem[   726] = 9'd31;    
		mem[   727] = 9'd28;    
		mem[   728] = 9'd66;    
		mem[   729] = 9'd28;    
		mem[   730] = 9'd30;    
		mem[   731] = 9'd62;    
		mem[   732] = 9'd31;    
		mem[   733] = 9'd29;    
		mem[   734] = 9'd65;    
		mem[   735] = 9'd28;    
		mem[   736] = 9'd29;    
		mem[   737] = 9'd63;    
		mem[   738] = 9'd31;    
		mem[   739] = 9'd29;    
		mem[   740] = 9'd36;    
		mem[   741] = 9'd29;    
		mem[   742] = 9'd28;    
		mem[   743] = 9'd30;    
		mem[   744] = 9'd62;    
		mem[   745] = 9'd31;    
		mem[   746] = 9'd29;    
		mem[   747] = 9'd35;    
		mem[   748] = 9'd30;    
		mem[   749] = 9'd29;    
		mem[   750] = 9'd29;    
		mem[   751] = 9'd62;    
		mem[   752] = 9'd31;    
		mem[   753] = 9'd29;    
		mem[   754] = 9'd35;    
		mem[   755] = 9'd30;    
		mem[   756] = 9'd29;    
		mem[   757] = 9'd29;    
		mem[   758] = 9'd35;    
		mem[   759] = 9'd28;    
		mem[   760] = 9'd31;    
		mem[   761] = 9'd29;    
		mem[   762] = 9'd34;    
		mem[   763] = 9'd29;    
		mem[   764] = 9'd30;    
		mem[   765] = 9'd17;    
		mem[   766] = 9'd13;    
		mem[   767] = 9'd62;    
		mem[   768] = 9'd31;    
		mem[   769] = 9'd17;    
		mem[   770] = 9'd12;    
		mem[   771] = 9'd32;    
		mem[   772] = 9'd30;    
		mem[   773] = 9'd32;    
		mem[   774] = 9'd30;    
		mem[   775] = 9'd31;    
		mem[   776] = 9'd30;    
		mem[   777] = 9'd31;    
		mem[   778] = 9'd30;    
		mem[   779] = 9'd32;    
		mem[   780] = 9'd30;    
		mem[   781] = 9'd31;    
		mem[   782] = 9'd30;    
		mem[   783] = 9'd31;    
		mem[   784] = 9'd30;    
		mem[   785] = 9'd31;    
		mem[   786] = 9'd30;    
		mem[   787] = 9'd32;    
		mem[   788] = 9'd29;    
		mem[   789] = 9'd32;    
		mem[   790] = 9'd30;    
		mem[   791] = 9'd31;    
		mem[   792] = 9'd30;    
		mem[   793] = 9'd31;    
		mem[   794] = 9'd30;    
		mem[   795] = 9'd32;    
		mem[   796] = 9'd32;    
		mem[   797] = 9'd33;    
		mem[   798] = 9'd32;    
		mem[   799] = 9'd33;    
		mem[   800] = 9'd32;    
		mem[   801] = 9'd33;    
		mem[   802] = 9'd32;    
		mem[   803] = 9'd33;    
		mem[   804] = 9'd32;    
		mem[   805] = 9'd33;    
		mem[   806] = 9'd32;    
		mem[   807] = 9'd33;    
		mem[   808] = 9'd32;    
		mem[   809] = 9'd33;    
		mem[   810] = 9'd32;    
		mem[   811] = 9'd33;    
		mem[   812] = 9'd32;    
		mem[   813] = 9'd33;    
		mem[   814] = 9'd32;    
		mem[   815] = 9'd33;    
		mem[   816] = 9'd32;    
		mem[   817] = 9'd33;    
		mem[   818] = 9'd30;    
		mem[   819] = 9'd31;    
		mem[   820] = 9'd30;    
		mem[   821] = 9'd32;    
		mem[   822] = 9'd29;    
		mem[   823] = 9'd32;    
		mem[   824] = 9'd30;    
		mem[   825] = 9'd31;    
		mem[   826] = 9'd30;    
		mem[   827] = 9'd31;    
		mem[   828] = 9'd30;    
		mem[   829] = 9'd31;    
		mem[   830] = 9'd30;    
		mem[   831] = 9'd32;    
		mem[   832] = 9'd30;    
		mem[   833] = 9'd31;    
		mem[   834] = 9'd30;    
		mem[   835] = 9'd31;    
		mem[   836] = 9'd30;    
		mem[   837] = 9'd32;    
		mem[   838] = 9'd30;    
		mem[   839] = 9'd31;    
		mem[   840] = 9'd30;    
		mem[   841] = 9'd64;    
		mem[   842] = 9'd27;    
		mem[   843] = 9'd92;    
		mem[   844] = 9'd31;    
		mem[   845] = 9'd94;    
		mem[   846] = 9'd28;    
		mem[   847] = 9'd92;    
		mem[   848] = 9'd31;    
		mem[   849] = 9'd94;    
		mem[   850] = 9'd28;    
		mem[   851] = 9'd92;    
		mem[   852] = 9'd31;    
		mem[   853] = 9'd94;    
		mem[   854] = 9'd29;    
		mem[   855] = 9'd29;    
		mem[   856] = 9'd63;    
		mem[   857] = 9'd30;    
		mem[   858] = 9'd94;    
		mem[   859] = 9'd29;    
		mem[   860] = 9'd29;    
		mem[   861] = 9'd63;    
		mem[   862] = 9'd30;    
		mem[   863] = 9'd29;    
		mem[   864] = 9'd65;    
		mem[   865] = 9'd29;    
		mem[   866] = 9'd29;    
		mem[   867] = 9'd63;    
		mem[   868] = 9'd31;    
		mem[   869] = 9'd28;    
		mem[   870] = 9'd63;    
		mem[   871] = 9'd31;    
		mem[   872] = 9'd31;    
		mem[   873] = 9'd31;    
		mem[   874] = 9'd30;    
		mem[   875] = 9'd32;    
		mem[   876] = 9'd30;    
		mem[   877] = 9'd31;    
		mem[   878] = 9'd30;    
		mem[   879] = 9'd31;    
		mem[   880] = 9'd30;    
		mem[   881] = 9'd32;    
		mem[   882] = 9'd29;    
		mem[   883] = 9'd32;    
		mem[   884] = 9'd30;    
		mem[   885] = 9'd31;    
		mem[   886] = 9'd30;    
		mem[   887] = 9'd31;    
		mem[   888] = 9'd30;    
		mem[   889] = 9'd32;    
		mem[   890] = 9'd29;    
		mem[   891] = 9'd32;    
		mem[   892] = 9'd30;    
		mem[   893] = 9'd67;    
		mem[   894] = 9'd63;    
		mem[   895] = 9'd48;    
		mem[   896] = 9'd19;    
		mem[   897] = 9'd62;    
		mem[   898] = 9'd65;    
		mem[   899] = 9'd67;    
		mem[   900] = 9'd30;    
		mem[   901] = 9'd32;    
		mem[   902] = 9'd67;    
		mem[   903] = 9'd62;    
		mem[   904] = 9'd69;    
		mem[   905] = 9'd49;    
		mem[   906] = 9'd78;    
		mem[   907] = 9'd30;    
		mem[   908] = 9'd15;    
		mem[   909] = 9'd77;    
		mem[   910] = 9'd36;    
		mem[   911] = 9'd11;    
		mem[   912] = 9'd11;    
		mem[   913] = 9'd66;    
		mem[   914] = 9'd30;    
		mem[   915] = 9'd14;    
		mem[   916] = 9'd77;    
		mem[   917] = 9'd36;    
		mem[   918] = 9'd11;    
		mem[   919] = 9'd11;    
		mem[   920] = 9'd66;    
		mem[   921] = 9'd30;    
		mem[   922] = 9'd14;    
		mem[   923] = 9'd12;    
		mem[   924] = 9'd65;    
		mem[   925] = 9'd36;    
		mem[   926] = 9'd11;    
		mem[   927] = 9'd11;    
		mem[   928] = 9'd65;    
		mem[   929] = 9'd31;    
		mem[   930] = 9'd15;    
		mem[   931] = 9'd12;    
		mem[   932] = 9'd64;    
		mem[   933] = 9'd36;    
		mem[   934] = 9'd23;    
		mem[   935] = 9'd65;    
		mem[   936] = 9'd30;    
		mem[   937] = 9'd15;    
		mem[   938] = 9'd12;    
		mem[   939] = 9'd36;    
		mem[   940] = 9'd28;    
		mem[   941] = 9'd36;    
		mem[   942] = 9'd23;    
		mem[   943] = 9'd64;    
		mem[   944] = 9'd14;    
		mem[   945] = 9'd17;    
		mem[   946] = 9'd15;    
		mem[   947] = 9'd12;    
		mem[   948] = 9'd36;    
		mem[   949] = 9'd28;    
		mem[   950] = 9'd36;    
		mem[   951] = 9'd23;    
		mem[   952] = 9'd64;    
		mem[   953] = 9'd31;    
		mem[   954] = 9'd16;    
		mem[   955] = 9'd11;    
		mem[   956] = 9'd36;    
		mem[   957] = 9'd28;    
		mem[   958] = 9'd36;    
		mem[   959] = 9'd23;    
		mem[   960] = 9'd31;    
		mem[   961] = 9'd34;    
		mem[   962] = 9'd30;    
		mem[   963] = 9'd27;    
		mem[   964] = 9'd35;    
		mem[   965] = 9'd29;    
		mem[   966] = 9'd33;    
		mem[   967] = 9'd27;    
		mem[   968] = 9'd31;    
		mem[   969] = 9'd32;    
		mem[   970] = 9'd31;    
		mem[   971] = 9'd28;    
		mem[   972] = 9'd34;    
		mem[   973] = 9'd29;    
		mem[   974] = 9'd33;    
		mem[   975] = 9'd26;    
		mem[   976] = 9'd62;    
		mem[   977] = 9'd31;    
		mem[   978] = 9'd31;    
		mem[   979] = 9'd31;    
		mem[   980] = 9'd30;    
		mem[   981] = 9'd32;    
		mem[   982] = 9'd30;    
		mem[   983] = 9'd31;    
		mem[   984] = 9'd30;    
		mem[   985] = 9'd32;    
		mem[   986] = 9'd30;    
		mem[   987] = 9'd31;    
		mem[   988] = 9'd30;    
		mem[   989] = 9'd31;    
		mem[   990] = 9'd30;    
		mem[   991] = 9'd31;    
		mem[   992] = 9'd30;    
		mem[   993] = 9'd31;    
		mem[   994] = 9'd30;    
		mem[   995] = 9'd32;    
		mem[   996] = 9'd30;    
		mem[   997] = 9'd31;    
		mem[   998] = 9'd33;    
		mem[   999] = 9'd39;    
		mem[  1000] = 9'd38;    
		mem[  1001] = 9'd40;    
		mem[  1002] = 9'd38;    
		mem[  1003] = 9'd40;    
		mem[  1004] = 9'd38;    
		mem[  1005] = 9'd39;    
		mem[  1006] = 9'd38;    
		mem[  1007] = 9'd40;    
		mem[  1008] = 9'd38;    
		mem[  1009] = 9'd39;    
		mem[  1010] = 9'd39;    
		mem[  1011] = 9'd39;    
		mem[  1012] = 9'd38;    
		mem[  1013] = 9'd40;    
		mem[  1014] = 9'd38;    
		mem[  1015] = 9'd40;    
		mem[  1016] = 9'd38;    
		mem[  1017] = 9'd38;    
		mem[  1018] = 9'd36;    
		mem[  1019] = 9'd37;    
		mem[  1020] = 9'd36;    
		mem[  1021] = 9'd37;    
		mem[  1022] = 9'd36;    
		mem[  1023] = 9'd37;    
		mem[  1024] = 9'd36;    
		mem[  1025] = 9'd38;    
		mem[  1026] = 9'd36;    
		mem[  1027] = 9'd37;    
		mem[  1028] = 9'd36;    
		mem[  1029] = 9'd37;    
		mem[  1030] = 9'd36;    
		mem[  1031] = 9'd37;    
		mem[  1032] = 9'd36;    
		mem[  1033] = 9'd37;    
		mem[  1034] = 9'd36;    
		mem[  1035] = 9'd38;    
		mem[  1036] = 9'd35;    
		mem[  1037] = 9'd37;    
		mem[  1038] = 9'd76;    
		mem[  1039] = 9'd102;    
		mem[  1040] = 9'd22;    
		mem[  1041] = 9'd55;    
		mem[  1042] = 9'd74;    
		mem[  1043] = 9'd75;    
		mem[  1044] = 9'd41;    
		mem[  1045] = 9'd106;    
		mem[  1046] = 9'd72;    
		mem[  1047] = 9'd37;    
		mem[  1048] = 9'd35;    
		mem[  1049] = 9'd83;    
		mem[  1050] = 9'd19;    
		mem[  1051] = 9'd19;    
		mem[  1052] = 9'd40;    
		mem[  1053] = 9'd46;    
		mem[  1054] = 9'd37;    
		mem[  1055] = 9'd85;    
		mem[  1056] = 9'd20;    
		mem[  1057] = 9'd18;    
		mem[  1058] = 9'd40;    
		mem[  1059] = 9'd46;    
		mem[  1060] = 9'd37;    
		mem[  1061] = 9'd85;    
		mem[  1062] = 9'd18;    
		mem[  1063] = 9'd20;    
		mem[  1064] = 9'd40;    
		mem[  1065] = 9'd46;    
		mem[  1066] = 9'd37;    
		mem[  1067] = 9'd41;    
		mem[  1068] = 9'd41;    
		mem[  1069] = 9'd41;    
		mem[  1070] = 9'd41;    
		mem[  1071] = 9'd41;    
		mem[  1072] = 9'd41;    
		mem[  1073] = 9'd41;    
		mem[  1074] = 9'd41;    
		mem[  1075] = 9'd41;    
		mem[  1076] = 9'd40;    
		mem[  1077] = 9'd42;    
		mem[  1078] = 9'd40;    
		mem[  1079] = 9'd42;    
		mem[  1080] = 9'd40;    
		mem[  1081] = 9'd42;    
		mem[  1082] = 9'd40;    
		mem[  1083] = 9'd42;    
		mem[  1084] = 9'd38;    
		mem[  1085] = 9'd64;    
		mem[  1086] = 9'd57;    
		mem[  1087] = 9'd66;    
		mem[  1088] = 9'd57;    
		mem[  1089] = 9'd65;    
		mem[  1090] = 9'd57;    
		mem[  1091] = 9'd66;    
		mem[  1092] = 9'd57;    
		mem[  1093] = 9'd65;    
		mem[  1094] = 9'd58;    
		mem[  1095] = 9'd65;    
		mem[  1096] = 9'd58;    
		mem[  1097] = 9'd64;    
		mem[  1098] = 9'd58;    
		mem[  1099] = 9'd65;    
		mem[  1100] = 9'd58;    
		mem[  1101] = 9'd64;    
		mem[  1102] = 9'd58;    
		mem[  1103] = 9'd65;    
		mem[  1104] = 9'd58;    
		mem[  1105] = 9'd64;    
		mem[  1106] = 9'd58;    
		mem[  1107] = 9'd65;    
		mem[  1108] = 9'd24;    
		mem[  1109] = 9'd36;    
		mem[  1110] = 9'd111;    
		mem[  1111] = 9'd91;    
		mem[  1112] = 9'd31;    
		mem[  1113] = 9'd121;    
		mem[  1114] = 9'd93;    
		mem[  1115] = 9'd31;    
		mem[  1116] = 9'd122;    
		mem[  1117] = 9'd92;    
		mem[  1118] = 9'd35;    
		mem[  1119] = 9'd62;    
		mem[  1120] = 9'd34;    
		mem[  1121] = 9'd27;    
		mem[  1122] = 9'd63;    
		mem[  1123] = 9'd29;    
		mem[  1124] = 9'd31;    
		mem[  1125] = 9'd62;    
		mem[  1126] = 9'd60;    
		mem[  1127] = 9'd63;    
		mem[  1128] = 9'd30;    
		mem[  1129] = 9'd30;    
		mem[  1130] = 9'd62;    
		mem[  1131] = 9'd34;    
		mem[  1132] = 9'd26;    
		mem[  1133] = 9'd63;    
		mem[  1134] = 9'd30;    
		mem[  1135] = 9'd28;    
		mem[  1136] = 9'd62;    
		mem[  1137] = 9'd31;    
		mem[  1138] = 9'd31;    
		mem[  1139] = 9'd32;    
		mem[  1140] = 9'd30;    
		mem[  1141] = 9'd31;    
		mem[  1142] = 9'd30;    
		mem[  1143] = 9'd32;    
		mem[  1144] = 9'd30;    
		mem[  1145] = 9'd31;    
		mem[  1146] = 9'd30;    
		mem[  1147] = 9'd32;    
		mem[  1148] = 9'd29;    
		mem[  1149] = 9'd32;    
		mem[  1150] = 9'd29;    
		mem[  1151] = 9'd32;    
		mem[  1152] = 9'd30;    
		mem[  1153] = 9'd31;    
		mem[  1154] = 9'd30;    
		mem[  1155] = 9'd31;    
		mem[  1156] = 9'd30;    
		mem[  1157] = 9'd32;    
		mem[  1158] = 9'd29;    
		mem[  1159] = 9'd32;    
		mem[  1160] = 9'd30;    
		mem[  1161] = 9'd31;    
		mem[  1162] = 9'd30;    
		mem[  1163] = 9'd31;    
		mem[  1164] = 9'd30;    
		mem[  1165] = 9'd31;    
		mem[  1166] = 9'd30;    
		mem[  1167] = 9'd32;    
		mem[  1168] = 9'd30;    
		mem[  1169] = 9'd31;    
		mem[  1170] = 9'd30;    
		mem[  1171] = 9'd31;    
		mem[  1172] = 9'd30;    
		mem[  1173] = 9'd31;    
		mem[  1174] = 9'd30;    
		mem[  1175] = 9'd32;    
		mem[  1176] = 9'd30;    
		mem[  1177] = 9'd31;    
		mem[  1178] = 9'd30;    
		mem[  1179] = 9'd31;    
		mem[  1180] = 9'd30;    
		mem[  1181] = 9'd31;    
		mem[  1182] = 9'd30;    
		mem[  1183] = 9'd31;    
		mem[  1184] = 9'd31;    
		mem[  1185] = 9'd31;    
		mem[  1186] = 9'd30;    
		mem[  1187] = 9'd31;    
		mem[  1188] = 9'd30;    
		mem[  1189] = 9'd31;    
		mem[  1190] = 9'd30;    
		mem[  1191] = 9'd32;    
		mem[  1192] = 9'd30;    
		mem[  1193] = 9'd31;    
		mem[  1194] = 9'd30;    
		mem[  1195] = 9'd31;    
		mem[  1196] = 9'd30;    
		mem[  1197] = 9'd31;    
		mem[  1198] = 9'd31;    
		mem[  1199] = 9'd31;    
		mem[  1200] = 9'd30;    
		mem[  1201] = 9'd31;    
		mem[  1202] = 9'd30;    
		mem[  1203] = 9'd31;    
		mem[  1204] = 9'd30;    
		mem[  1205] = 9'd72;    
		mem[  1206] = 9'd81;    
		mem[  1207] = 9'd79;    
		mem[  1208] = 9'd57;    
		mem[  1209] = 9'd58;    
		mem[  1210] = 9'd39;    
		mem[  1211] = 9'd78;    
		mem[  1212] = 9'd35;    
		mem[  1213] = 9'd38;    
		mem[  1214] = 9'd83;    
		mem[  1215] = 9'd35;    
		mem[  1216] = 9'd39;    
		mem[  1217] = 9'd43;    
		mem[  1218] = 9'd35;    
		mem[  1219] = 9'd74;    
		mem[  1220] = 9'd39;    
		mem[  1221] = 9'd17;    
		mem[  1222] = 9'd88;    
		mem[  1223] = 9'd35;    
		mem[  1224] = 9'd37;    
		mem[  1225] = 9'd75;    
		mem[  1226] = 9'd76;    
		mem[  1227] = 9'd68;    
		mem[  1228] = 9'd38;    
		mem[  1229] = 9'd40;    
		mem[  1230] = 9'd32;    
		mem[  1231] = 9'd38;    
		mem[  1232] = 9'd41;    
		mem[  1233] = 9'd34;    
		mem[  1234] = 9'd38;    
		mem[  1235] = 9'd34;    
		mem[  1236] = 9'd37;    
		mem[  1237] = 9'd36;    
		mem[  1238] = 9'd37;    
		mem[  1239] = 9'd36;    
		mem[  1240] = 9'd37;    
		mem[  1241] = 9'd36;    
		mem[  1242] = 9'd37;    
		mem[  1243] = 9'd36;    
		mem[  1244] = 9'd37;    
		mem[  1245] = 9'd37;    
		mem[  1246] = 9'd36;    
		mem[  1247] = 9'd37;    
		mem[  1248] = 9'd37;    
		mem[  1249] = 9'd36;    
		mem[  1250] = 9'd37;    
		mem[  1251] = 9'd36;    
		mem[  1252] = 9'd37;    
		mem[  1253] = 9'd35;    
		mem[  1254] = 9'd77;    
		mem[  1255] = 9'd74;    
		mem[  1256] = 9'd40;    
		mem[  1257] = 9'd103;    
		mem[  1258] = 9'd73;    
		mem[  1259] = 9'd19;    
		mem[  1260] = 9'd55;    
		mem[  1261] = 9'd39;    
		mem[  1262] = 9'd16;    
		mem[  1263] = 9'd61;    
		mem[  1264] = 9'd7;    
		mem[  1265] = 9'd23;    
		mem[  1266] = 9'd76;    
		mem[  1267] = 9'd73;    
		mem[  1268] = 9'd14;    
		mem[  1269] = 9'd20;    
		mem[  1270] = 9'd20;    
		mem[  1271] = 9'd13;    
		mem[  1272] = 9'd76;    
		mem[  1273] = 9'd73;    
		mem[  1274] = 9'd22;    
		mem[  1275] = 9'd52;    
		mem[  1276] = 9'd40;    
		mem[  1277] = 9'd16;    
		mem[  1278] = 9'd58;    
		mem[  1279] = 9'd12;    
		mem[  1280] = 9'd20;    
		mem[  1281] = 9'd76;    
		mem[  1282] = 9'd73;    
		mem[  1283] = 9'd14;    
		mem[  1284] = 9'd41;    
		mem[  1285] = 9'd13;    
		mem[  1286] = 9'd77;    
		mem[  1287] = 9'd38;    
		mem[  1288] = 9'd35;    
		mem[  1289] = 9'd37;    
		mem[  1290] = 9'd35;    
		mem[  1291] = 9'd37;    
		mem[  1292] = 9'd36;    
		mem[  1293] = 9'd37;    
		mem[  1294] = 9'd36;    
		mem[  1295] = 9'd39;    
		mem[  1296] = 9'd33;    
		mem[  1297] = 9'd72;    
		mem[  1298] = 9'd78;    
		mem[  1299] = 9'd34;    
		mem[  1300] = 9'd38;    
		mem[  1301] = 9'd34;    
		mem[  1302] = 9'd25;    
		mem[  1303] = 9'd87;    
		mem[  1304] = 9'd72;    
		mem[  1305] = 9'd19;    
		mem[  1306] = 9'd56;    
		mem[  1307] = 9'd37;    
		mem[  1308] = 9'd35;    
		mem[  1309] = 9'd37;    
		mem[  1310] = 9'd34;    
		mem[  1311] = 9'd76;    
		mem[  1312] = 9'd73;    
		mem[  1313] = 9'd74;    
		mem[  1314] = 9'd38;    
		mem[  1315] = 9'd32;    
		mem[  1316] = 9'd40;    
		mem[  1317] = 9'd33;    
		mem[  1318] = 9'd40;    
		mem[  1319] = 9'd36;    
		mem[  1320] = 9'd73;    
		mem[  1321] = 9'd33;    
		mem[  1322] = 9'd40;    
		mem[  1323] = 9'd39;    
		mem[  1324] = 9'd17;    
		mem[  1325] = 9'd15;    
		mem[  1326] = 9'd42;    
		mem[  1327] = 9'd32;    
		mem[  1328] = 9'd59;    
		mem[  1329] = 9'd14;    
		mem[  1330] = 9'd37;    
		mem[  1331] = 9'd37;    
		mem[  1332] = 9'd37;    
		mem[  1333] = 9'd36;    
		mem[  1334] = 9'd38;    
		mem[  1335] = 9'd36;    
		mem[  1336] = 9'd37;    
		mem[  1337] = 9'd36;    
		mem[  1338] = 9'd75;    
		mem[  1339] = 9'd71;    
		mem[  1340] = 9'd20;    
		mem[  1341] = 9'd56;    
		mem[  1342] = 9'd34;    
		mem[  1343] = 9'd38;    
		mem[  1344] = 9'd30;    
		mem[  1345] = 9'd25;    
		mem[  1346] = 9'd87;    
		mem[  1347] = 9'd62;    
		mem[  1348] = 9'd16;    
		mem[  1349] = 9'd73;    
		mem[  1350] = 9'd73;    
		mem[  1351] = 9'd34;    
		mem[  1352] = 9'd36;    
		mem[  1353] = 9'd41;    
		mem[  1354] = 9'd70;    
		mem[  1355] = 9'd23;    
		mem[  1356] = 9'd87;    
		mem[  1357] = 9'd68;    
		mem[  1358] = 9'd22;    
		mem[  1359] = 9'd84;    
		mem[  1360] = 9'd68;    
		mem[  1361] = 9'd22;    
		mem[  1362] = 9'd85;    
		mem[  1363] = 9'd67;    
		mem[  1364] = 9'd23;    
		mem[  1365] = 9'd84;    
		mem[  1366] = 9'd430;    
		mem[  1367] = 9'd21;    
		mem[  1368] = 9'd80;    
		mem[  1369] = 9'd61;    
		mem[  1370] = 9'd19;    
		mem[  1371] = 9'd81;    
		mem[  1372] = 9'd61;    
		mem[  1373] = 9'd22;    
		mem[  1374] = 9'd81;    
		mem[  1375] = 9'd61;    
		mem[  1376] = 9'd21;    
		mem[  1377] = 9'd82;    
		mem[  1378] = 9'd62;    
		mem[  1379] = 9'd21;    
		mem[  1380] = 9'd80;    
		mem[  1381] = 9'd62;    
		mem[  1382] = 9'd22;    
		mem[  1383] = 9'd80;    
		mem[  1384] = 9'd64;    
		mem[  1385] = 9'd20;    
		mem[  1386] = 9'd80;    
		mem[  1387] = 9'd64;    
		mem[  1388] = 9'd20;    
		mem[  1389] = 9'd80;    
		mem[  1390] = 9'd62;    
		mem[  1391] = 9'd22;    
		mem[  1392] = 9'd250;    
		mem[  1393] = 9'd197;    
		mem[  1394] = 9'd97;    
		mem[  1395] = 9'd33;    
		mem[  1396] = 9'd100;    
		mem[  1397] = 9'd63;    
		mem[  1398] = 9'd52;    
		mem[  1399] = 9'd13;    
		mem[  1400] = 9'd64;    
		mem[  1401] = 9'd66;    
		mem[  1402] = 9'd67;    
		mem[  1403] = 9'd30;    
		mem[  1404] = 9'd33;    
		mem[  1405] = 9'd66;    
		mem[  1406] = 9'd61;    
		mem[  1407] = 9'd65;    
		mem[  1408] = 9'd25;    
		mem[  1409] = 9'd33;    
		mem[  1410] = 9'd63;    
		mem[  1411] = 9'd59;    
		mem[  1412] = 9'd65;    
		mem[  1413] = 9'd26;    
		mem[  1414] = 9'd32;    
		mem[  1415] = 9'd63;    
		mem[  1416] = 9'd59;    
		mem[  1417] = 9'd65;    
		mem[  1418] = 9'd26;    
		mem[  1419] = 9'd32;    
		mem[  1420] = 9'd63;    
		mem[  1421] = 9'd59;    
		mem[  1422] = 9'd64;    
		mem[  1423] = 9'd27;    
		mem[  1424] = 9'd32;    
		mem[  1425] = 9'd63;    
		mem[  1426] = 9'd59;    
		mem[  1427] = 9'd65;    
		mem[  1428] = 9'd26;    
		mem[  1429] = 9'd32;    
		mem[  1430] = 9'd63;    
		mem[  1431] = 9'd59;    
		mem[  1432] = 9'd64;    
		mem[  1433] = 9'd27;    
		mem[  1434] = 9'd32;    
		mem[  1435] = 9'd63;    
		mem[  1436] = 9'd60;    
		mem[  1437] = 9'd63;    
		mem[  1438] = 9'd27;    
		mem[  1439] = 9'd32;    
		mem[  1440] = 9'd63;    
		mem[  1441] = 9'd34;    
		mem[  1442] = 9'd26;    
		mem[  1443] = 9'd64;    
		mem[  1444] = 9'd27;    
		mem[  1445] = 9'd31;    
		mem[  1446] = 9'd63;    
		mem[  1447] = 9'd33;    
		mem[  1448] = 9'd27;    
		mem[  1449] = 9'd63;    
		mem[  1450] = 9'd28;    
		mem[  1451] = 9'd32;    
		mem[  1452] = 9'd62;    
		mem[  1453] = 9'd62;    
		mem[  1454] = 9'd32;    
		mem[  1455] = 9'd28;    
		mem[  1456] = 9'd32;    
		mem[  1457] = 9'd29;    
		mem[  1458] = 9'd31;    
		mem[  1459] = 9'd30;    
		mem[  1460] = 9'd31;    
		mem[  1461] = 9'd30;    
		mem[  1462] = 9'd31;    
		mem[  1463] = 9'd31;    
		mem[  1464] = 9'd30;    
		mem[  1465] = 9'd31;    
		mem[  1466] = 9'd30;    
		mem[  1467] = 9'd31;    
		mem[  1468] = 9'd31;    
		mem[  1469] = 9'd31;    
		mem[  1470] = 9'd30;    
		mem[  1471] = 9'd31;    
		mem[  1472] = 9'd31;    
		mem[  1473] = 9'd30;    
		mem[  1474] = 9'd31;    
		mem[  1475] = 9'd31;    
		mem[  1476] = 9'd32;    
		mem[  1477] = 9'd32;    
		mem[  1478] = 9'd33;    
		mem[  1479] = 9'd32;    
		mem[  1480] = 9'd33;    
		mem[  1481] = 9'd32;    
		mem[  1482] = 9'd33;    
		mem[  1483] = 9'd32;    
		mem[  1484] = 9'd33;    
		mem[  1485] = 9'd32;    
		mem[  1486] = 9'd33;    
		mem[  1487] = 9'd32;    
		mem[  1488] = 9'd33;    
		mem[  1489] = 9'd32;    
		mem[  1490] = 9'd33;    
		mem[  1491] = 9'd32;    
		mem[  1492] = 9'd33;    
		mem[  1493] = 9'd32;    
		mem[  1494] = 9'd33;    
		mem[  1495] = 9'd32;    
		mem[  1496] = 9'd33;    
		mem[  1497] = 9'd32;    
		mem[  1498] = 9'd33;    
		mem[  1499] = 9'd30;    
		mem[  1500] = 9'd31;    
		mem[  1501] = 9'd30;    
		mem[  1502] = 9'd31;    
		mem[  1503] = 9'd30;    
		mem[  1504] = 9'd31;    
		mem[  1505] = 9'd30;    
		mem[  1506] = 9'd31;    
		mem[  1507] = 9'd30;    
		mem[  1508] = 9'd31;    
		mem[  1509] = 9'd31;    
		mem[  1510] = 9'd31;    
		mem[  1511] = 9'd30;    
		mem[  1512] = 9'd31;    
		mem[  1513] = 9'd30;    
		mem[  1514] = 9'd31;    
		mem[  1515] = 9'd30;    
		mem[  1516] = 9'd32;    
		mem[  1517] = 9'd30;    
		mem[  1518] = 9'd31;    
		mem[  1519] = 9'd30;    
		mem[  1520] = 9'd31;    
		mem[  1521] = 9'd30;    
		mem[  1522] = 9'd32;    
		mem[  1523] = 9'd27;    
		mem[  1524] = 9'd66;    
		mem[  1525] = 9'd26;    
		mem[  1526] = 9'd32;    
		mem[  1527] = 9'd64;    
		mem[  1528] = 9'd58;    
		mem[  1529] = 9'd66;    
		mem[  1530] = 9'd12;    
		mem[  1531] = 9'd13;    
		mem[  1532] = 9'd32;    
		mem[  1533] = 9'd64;    
		mem[  1534] = 9'd59;    
		mem[  1535] = 9'd65;    
		mem[  1536] = 9'd11;    
		mem[  1537] = 9'd14;    
		mem[  1538] = 9'd32;    
		mem[  1539] = 9'd64;    
		mem[  1540] = 9'd59;    
		mem[  1541] = 9'd65;    
		mem[  1542] = 9'd25;    
		mem[  1543] = 9'd32;    
		mem[  1544] = 9'd64;    
		mem[  1545] = 9'd58;    
		mem[  1546] = 9'd65;    
		mem[  1547] = 9'd26;    
		mem[  1548] = 9'd32;    
		mem[  1549] = 9'd64;    
		mem[  1550] = 9'd59;    
		mem[  1551] = 9'd64;    
		mem[  1552] = 9'd26;    
		mem[  1553] = 9'd33;    
		mem[  1554] = 9'd63;    
		mem[  1555] = 9'd33;    
		mem[  1556] = 9'd28;    
		mem[  1557] = 9'd31;    
		mem[  1558] = 9'd30;    
		mem[  1559] = 9'd31;    
		mem[  1560] = 9'd30;    
		mem[  1561] = 9'd31;    
		mem[  1562] = 9'd30;    
		mem[  1563] = 9'd31;    
		mem[  1564] = 9'd30;    
		mem[  1565] = 9'd31;    
		mem[  1566] = 9'd30;    
		mem[  1567] = 9'd31;    
		mem[  1568] = 9'd30;    
		mem[  1569] = 9'd31;    
		mem[  1570] = 9'd31;    
		mem[  1571] = 9'd31;    
		mem[  1572] = 9'd30;    
		mem[  1573] = 9'd31;    
		mem[  1574] = 9'd30;    
		mem[  1575] = 9'd31;    
		mem[  1576] = 9'd31;    
		mem[  1577] = 9'd31;    
		mem[  1578] = 9'd31;    
		mem[  1579] = 9'd34;    
		mem[  1580] = 9'd96;    
		mem[  1581] = 9'd36;    
		mem[  1582] = 9'd62;    
		mem[  1583] = 9'd34;    
		mem[  1584] = 9'd29;    
		mem[  1585] = 9'd97;    
		mem[  1586] = 9'd32;    
		mem[  1587] = 9'd32;    
		mem[  1588] = 9'd69;    
		mem[  1589] = 9'd63;    
		mem[  1590] = 9'd36;    
		mem[  1591] = 9'd13;    
		mem[  1592] = 9'd18;    
		mem[  1593] = 9'd62;    
		mem[  1594] = 9'd63;    
		mem[  1595] = 9'd62;    
		mem[  1596] = 9'd31;    
		mem[  1597] = 9'd31;    
		mem[  1598] = 9'd59;    
		mem[  1599] = 9'd62;    
		mem[  1600] = 9'd62;    
		mem[  1601] = 9'd31;    
		mem[  1602] = 9'd30;    
		mem[  1603] = 9'd60;    
		mem[  1604] = 9'd62;    
		mem[  1605] = 9'd62;    
		mem[  1606] = 9'd31;    
		mem[  1607] = 9'd31;    
		mem[  1608] = 9'd59;    
		mem[  1609] = 9'd62;    
		mem[  1610] = 9'd62;    
		mem[  1611] = 9'd31;    
		mem[  1612] = 9'd31;    
		mem[  1613] = 9'd59;    
		mem[  1614] = 9'd62;    
		mem[  1615] = 9'd62;    
		mem[  1616] = 9'd31;    
		mem[  1617] = 9'd31;    
		mem[  1618] = 9'd59;    
		mem[  1619] = 9'd62;    
		mem[  1620] = 9'd62;    
		mem[  1621] = 9'd31;    
		mem[  1622] = 9'd31;    
		mem[  1623] = 9'd59;    
		mem[  1624] = 9'd62;    
		mem[  1625] = 9'd62;    
		mem[  1626] = 9'd31;    
		mem[  1627] = 9'd31;    
		mem[  1628] = 9'd59;    
		mem[  1629] = 9'd62;    
		mem[  1630] = 9'd62;    
		mem[  1631] = 9'd31;    
		mem[  1632] = 9'd30;    
		mem[  1633] = 9'd60;    
		mem[  1634] = 9'd62;    
		mem[  1635] = 9'd62;    
		mem[  1636] = 9'd31;    
		mem[  1637] = 9'd31;    
		mem[  1638] = 9'd46;    
		mem[  1639] = 9'd12;    
		mem[  1640] = 9'd62;    
		mem[  1641] = 9'd31;    
		mem[  1642] = 9'd31;    
		mem[  1643] = 9'd31;    
		mem[  1644] = 9'd30;    
		mem[  1645] = 9'd32;    
		mem[  1646] = 9'd30;    
		mem[  1647] = 9'd31;    
		mem[  1648] = 9'd30;    
		mem[  1649] = 9'd32;    
		mem[  1650] = 9'd29;    
		mem[  1651] = 9'd32;    
		mem[  1652] = 9'd30;    
		mem[  1653] = 9'd31;    
		mem[  1654] = 9'd30;    
		mem[  1655] = 9'd31;    
		mem[  1656] = 9'd30;    
		mem[  1657] = 9'd32;    
		mem[  1658] = 9'd29;    
		mem[  1659] = 9'd32;    
		mem[  1660] = 9'd30;    
		mem[  1661] = 9'd31;    
		mem[  1662] = 9'd36;    
		mem[  1663] = 9'd39;    
		mem[  1664] = 9'd38;    
		mem[  1665] = 9'd40;    
		mem[  1666] = 9'd38;    
		mem[  1667] = 9'd40;    
		mem[  1668] = 9'd38;    
		mem[  1669] = 9'd39;    
		mem[  1670] = 9'd38;    
		mem[  1671] = 9'd40;    
		mem[  1672] = 9'd38;    
		mem[  1673] = 9'd40;    
		mem[  1674] = 9'd38;    
		mem[  1675] = 9'd39;    
		mem[  1676] = 9'd38;    
		mem[  1677] = 9'd40;    
		mem[  1678] = 9'd38;    
		mem[  1679] = 9'd39;    
		mem[  1680] = 9'd39;    
		mem[  1681] = 9'd37;    
		mem[  1682] = 9'd36;    
		mem[  1683] = 9'd37;    
		mem[  1684] = 9'd36;    
		mem[  1685] = 9'd37;    
		mem[  1686] = 9'd36;    
		mem[  1687] = 9'd38;    
		mem[  1688] = 9'd35;    
		mem[  1689] = 9'd38;    
		mem[  1690] = 9'd36;    
		mem[  1691] = 9'd37;    
		mem[  1692] = 9'd36;    
		mem[  1693] = 9'd37;    
		mem[  1694] = 9'd36;    
		mem[  1695] = 9'd37;    
		mem[  1696] = 9'd36;    
		mem[  1697] = 9'd37;    
		mem[  1698] = 9'd36;    
		mem[  1699] = 9'd37;    
		mem[  1700] = 9'd36;    
		mem[  1701] = 9'd75;    
		mem[  1702] = 9'd75;    
		mem[  1703] = 9'd14;    
		mem[  1704] = 9'd14;    
		mem[  1705] = 9'd39;    
		mem[  1706] = 9'd79;    
		mem[  1707] = 9'd32;    
		mem[  1708] = 9'd80;    
		mem[  1709] = 9'd15;    
		mem[  1710] = 9'd18;    
		mem[  1711] = 9'd72;    
		mem[  1712] = 9'd70;    
		mem[  1713] = 9'd77;    
		mem[  1714] = 9'd35;    
		mem[  1715] = 9'd119;    
		mem[  1716] = 9'd84;    
		mem[  1717] = 9'd40;    
		mem[  1718] = 9'd122;    
		mem[  1719] = 9'd83;    
		mem[  1720] = 9'd41;    
		mem[  1721] = 9'd38;    
		mem[  1722] = 9'd84;    
		mem[  1723] = 9'd83;    
		mem[  1724] = 9'd40;    
		mem[  1725] = 9'd122;    
		mem[  1726] = 9'd42;    
		mem[  1727] = 9'd40;    
		mem[  1728] = 9'd43;    
		mem[  1729] = 9'd40;    
		mem[  1730] = 9'd42;    
		mem[  1731] = 9'd40;    
		mem[  1732] = 9'd42;    
		mem[  1733] = 9'd40;    
		mem[  1734] = 9'd42;    
		mem[  1735] = 9'd39;    
		mem[  1736] = 9'd42;    
		mem[  1737] = 9'd40;    
		mem[  1738] = 9'd42;    
		mem[  1739] = 9'd40;    
		mem[  1740] = 9'd42;    
		mem[  1741] = 9'd35;    
		mem[  1742] = 9'd64;    
		mem[  1743] = 9'd58;    
		mem[  1744] = 9'd54;    
		mem[  1745] = 9'd22;    
		mem[  1746] = 9'd109;    
		mem[  1747] = 9'd60;    
		mem[  1748] = 9'd54;    
		mem[  1749] = 9'd22;    
		mem[  1750] = 9'd44;    
		mem[  1751] = 9'd65;    
		mem[  1752] = 9'd60;    
		mem[  1753] = 9'd54;    
		mem[  1754] = 9'd22;    
		mem[  1755] = 9'd45;    
		mem[  1756] = 9'd64;    
		mem[  1757] = 9'd60;    
		mem[  1758] = 9'd55;    
		mem[  1759] = 9'd21;    
		mem[  1760] = 9'd45;    
		mem[  1761] = 9'd65;    
		mem[  1762] = 9'd59;    
		mem[  1763] = 9'd58;    
		mem[  1764] = 9'd18;    
		mem[  1765] = 9'd45;    
		mem[  1766] = 9'd64;    
		mem[  1767] = 9'd60;    
		mem[  1768] = 9'd58;    
		mem[  1769] = 9'd18;    
		mem[  1770] = 9'd123;    
		mem[  1771] = 9'd93;    
		mem[  1772] = 9'd32;    
		mem[  1773] = 9'd121;    
		mem[  1774] = 9'd93;    
		mem[  1775] = 9'd32;    
		mem[  1776] = 9'd120;    
		mem[  1777] = 9'd93;    
		mem[  1778] = 9'd31;    
		mem[  1779] = 9'd37;    
		mem[  1780] = 9'd64;    
		mem[  1781] = 9'd28;    
		mem[  1782] = 9'd30;    
		mem[  1783] = 9'd61;    
		mem[  1784] = 9'd31;    
		mem[  1785] = 9'd30;    
		mem[  1786] = 9'd35;    
		mem[  1787] = 9'd29;    
		mem[  1788] = 9'd28;    
		mem[  1789] = 9'd31;    
		mem[  1790] = 9'd35;    
		mem[  1791] = 9'd27;    
		mem[  1792] = 9'd30;    
		mem[  1793] = 9'd19;    
		mem[  1794] = 9'd12;    
		mem[  1795] = 9'd34;    
		mem[  1796] = 9'd29;    
		mem[  1797] = 9'd29;    
		mem[  1798] = 9'd31;    
		mem[  1799] = 9'd35;    
		mem[  1800] = 9'd26;    
		mem[  1801] = 9'd32;    
		mem[  1802] = 9'd30;    
		mem[  1803] = 9'd31;    
		mem[  1804] = 9'd30;    
		mem[  1805] = 9'd31;    
		mem[  1806] = 9'd30;    
		mem[  1807] = 9'd31;    
		mem[  1808] = 9'd31;    
		mem[  1809] = 9'd31;    
		mem[  1810] = 9'd30;    
		mem[  1811] = 9'd31;    
		mem[  1812] = 9'd30;    
		mem[  1813] = 9'd31;    
		mem[  1814] = 9'd30;    
		mem[  1815] = 9'd31;    
		mem[  1816] = 9'd31;    
		mem[  1817] = 9'd31;    
		mem[  1818] = 9'd30;    
		mem[  1819] = 9'd31;    
		mem[  1820] = 9'd30;    
		mem[  1821] = 9'd31;    
		mem[  1822] = 9'd30;    
		mem[  1823] = 9'd32;    
		mem[  1824] = 9'd30;    
		mem[  1825] = 9'd31;    
		mem[  1826] = 9'd30;    
		mem[  1827] = 9'd31;    
		mem[  1828] = 9'd30;    
		mem[  1829] = 9'd32;    
		mem[  1830] = 9'd30;    
		mem[  1831] = 9'd31;    
		mem[  1832] = 9'd30;    
		mem[  1833] = 9'd31;    
		mem[  1834] = 9'd30;    
		mem[  1835] = 9'd31;    
		mem[  1836] = 9'd30;    
		mem[  1837] = 9'd31;    
		mem[  1838] = 9'd31;    
		mem[  1839] = 9'd31;    
		mem[  1840] = 9'd30;    
		mem[  1841] = 9'd31;    
		mem[  1842] = 9'd30;    
		mem[  1843] = 9'd31;    
		mem[  1844] = 9'd31;    
		mem[  1845] = 9'd31;    
		mem[  1846] = 9'd30;    
		mem[  1847] = 9'd31;    
		mem[  1848] = 9'd30;    
		mem[  1849] = 9'd31;    
		mem[  1850] = 9'd30;    
		mem[  1851] = 9'd32;    
		mem[  1852] = 9'd30;    
		mem[  1853] = 9'd31;    
		mem[  1854] = 9'd30;    
		mem[  1855] = 9'd31;    
		mem[  1856] = 9'd30;    
		mem[  1857] = 9'd31;    
		mem[  1858] = 9'd30;    
		mem[  1859] = 9'd32;    
		mem[  1860] = 9'd30;    
		mem[  1861] = 9'd30;    
		mem[  1862] = 9'd31;    
		mem[  1863] = 9'd31;    
		mem[  1864] = 9'd30;    
		mem[  1865] = 9'd31;    
		mem[  1866] = 9'd30;    
		mem[  1867] = 9'd32;    
		mem[  1868] = 9'd30;    
		mem[  1869] = 9'd31;    
		mem[  1870] = 9'd30;    
		mem[  1871] = 9'd31;    
		mem[  1872] = 9'd30;    
		mem[  1873] = 9'd55;    
		mem[  1874] = 9'd57;    
		mem[  1875] = 9'd52;    
		mem[  1876] = 9'd55;    
		mem[  1877] = 9'd29;    
		mem[  1878] = 9'd83;    
		mem[  1879] = 9'd50;    
		mem[  1880] = 9'd59;    
		mem[  1881] = 9'd14;    
		mem[  1882] = 9'd11;    
		mem[  1883] = 9'd28;    
		mem[  1884] = 9'd54;    
		mem[  1885] = 9'd56;    
		mem[  1886] = 9'd52;    
		mem[  1887] = 9'd56;    
		mem[  1888] = 9'd28;    
		mem[  1889] = 9'd78;    
		mem[  1890] = 9'd50;    
		mem[  1891] = 9'd53;    
		mem[  1892] = 9'd27;    
		mem[  1893] = 9'd12;    
		mem[  1894] = 9'd11;    
		mem[  1895] = 9'd12;    
		mem[  1896] = 9'd68;    
		mem[  1897] = 9'd26;    
		mem[  1898] = 9'd25;    
		mem[  1899] = 9'd12;    
		mem[  1900] = 9'd10;    
		mem[  1901] = 9'd56;    
		mem[  1902] = 9'd23;    
		mem[  1903] = 9'd27;    
		mem[  1904] = 9'd50;    
		mem[  1905] = 9'd54;    
		mem[  1906] = 9'd24;    
		mem[  1907] = 9'd79;    
		mem[  1908] = 9'd25;    
		mem[  1909] = 9'd25;    
		mem[  1910] = 9'd27;    
		mem[  1911] = 9'd25;    
		mem[  1912] = 9'd26;    
		mem[  1913] = 9'd26;    
		mem[  1914] = 9'd26;    
		mem[  1915] = 9'd25;    
		mem[  1916] = 9'd26;    
		mem[  1917] = 9'd26;    
		mem[  1918] = 9'd26;    
		mem[  1919] = 9'd25;    
		mem[  1920] = 9'd27;    
		mem[  1921] = 9'd25;    
		mem[  1922] = 9'd26;    
		mem[  1923] = 9'd26;    
		mem[  1924] = 9'd26;    
		mem[  1925] = 9'd25;    
		mem[  1926] = 9'd26;    
		mem[  1927] = 9'd26;    
		mem[  1928] = 9'd26;    
		mem[  1929] = 9'd26;    
		mem[  1930] = 9'd26;    
		mem[  1931] = 9'd25;    
		mem[  1932] = 9'd26;    
		mem[  1933] = 9'd26;    
		mem[  1934] = 9'd26;    
		mem[  1935] = 9'd26;    
		mem[  1936] = 9'd26;    
		mem[  1937] = 9'd24;    
		mem[  1938] = 9'd55;    
		mem[  1939] = 9'd28;    
		mem[  1940] = 9'd19;    
		mem[  1941] = 9'd55;    
		mem[  1942] = 9'd29;    
		mem[  1943] = 9'd10;    
		mem[  1944] = 9'd66;    
		mem[  1945] = 9'd23;    
		mem[  1946] = 9'd77;    
		mem[  1947] = 9'd26;    
		mem[  1948] = 9'd79;    
		mem[  1949] = 9'd50;    
		mem[  1950] = 9'd42;    
		mem[  1951] = 9'd10;    
		mem[  1952] = 9'd50;    
		mem[  1953] = 9'd54;    
		mem[  1954] = 9'd53;    
		mem[  1955] = 9'd24;    
		mem[  1956] = 9'd25;    
		mem[  1957] = 9'd52;    
		mem[  1958] = 9'd51;    
		mem[  1959] = 9'd54;    
		mem[  1960] = 9'd49;    
		mem[  1961] = 9'd54;    
		mem[  1962] = 9'd27;    
		mem[  1963] = 9'd12;    
		mem[  1964] = 9'd9;    
		mem[  1965] = 9'd55;    
		mem[  1966] = 9'd27;    
		mem[  1967] = 9'd21;    
		mem[  1968] = 9'd29;    
		mem[  1969] = 9'd27;    
		mem[  1970] = 9'd24;    
		mem[  1971] = 9'd24;    
		mem[  1972] = 9'd52;    
		mem[  1973] = 9'd26;    
		mem[  1974] = 9'd25;    
		mem[  1975] = 9'd56;    
		mem[  1976] = 9'd47;    
		mem[  1977] = 9'd26;    
		mem[  1978] = 9'd23;    
		mem[  1979] = 9'd25;    
		mem[  1980] = 9'd23;    
		mem[  1981] = 9'd25;    
		mem[  1982] = 9'd24;    
		mem[  1983] = 9'd24;    
		mem[  1984] = 9'd25;    
		mem[  1985] = 9'd24;    
		mem[  1986] = 9'd24;    
		mem[  1987] = 9'd25;    
		mem[  1988] = 9'd24;    
		mem[  1989] = 9'd99;    
		mem[  1990] = 9'd26;    
		mem[  1991] = 9'd74;    
		mem[  1992] = 9'd10;    
		mem[  1993] = 9'd11;    
		mem[  1994] = 9'd73;    
		mem[  1995] = 9'd25;    
		mem[  1996] = 9'd75;    
		mem[  1997] = 9'd44;    
		mem[  1998] = 9'd44;    
		mem[  1999] = 9'd15;    
		mem[  2000] = 9'd33;    
		mem[  2001] = 9'd49;    
		mem[  2002] = 9'd44;    
		mem[  2003] = 9'd44;    
		mem[  2004] = 9'd15;    
		mem[  2005] = 9'd33;    
		mem[  2006] = 9'd49;    
		mem[  2007] = 9'd44;    
		mem[  2008] = 9'd44;    
		mem[  2009] = 9'd15;    
		mem[  2010] = 9'd33;    
		mem[  2011] = 9'd49;    
		mem[  2012] = 9'd44;    
		mem[  2013] = 9'd44;    
		mem[  2014] = 9'd15;    
		mem[  2015] = 9'd33;    
		mem[  2016] = 9'd49;    
		mem[  2017] = 9'd44;    
		mem[  2018] = 9'd44;    
		mem[  2019] = 9'd14;    
		mem[  2020] = 9'd34;    
		mem[  2021] = 9'd49;    
		mem[  2022] = 9'd44;    
		mem[  2023] = 9'd44;    
		mem[  2024] = 9'd14;    
		mem[  2025] = 9'd34;    
		mem[  2026] = 9'd48;    
		mem[  2027] = 9'd24;    
		mem[  2028] = 9'd22;    
		mem[  2029] = 9'd24;    
		mem[  2030] = 9'd22;    
		mem[  2031] = 9'd23;    
		mem[  2032] = 9'd23;    
		mem[  2033] = 9'd23;    
		mem[  2034] = 9'd23;    
		mem[  2035] = 9'd23;    
		mem[  2036] = 9'd23;    
		mem[  2037] = 9'd23;    
		mem[  2038] = 9'd23;    
		mem[  2039] = 9'd24;    
		mem[  2040] = 9'd23;    
		mem[  2041] = 9'd25;    
		mem[  2042] = 9'd21;    
		mem[  2043] = 9'd47;    
		mem[  2044] = 9'd23;    
		mem[  2045] = 9'd22;    
		mem[  2046] = 9'd47;    
		mem[  2047] = 9'd45;    
		mem[  2048] = 9'd49;    
		mem[  2049] = 9'd43;    
		mem[  2050] = 9'd50;    
		mem[  2051] = 9'd23;    
		mem[  2052] = 9'd11;    
		mem[  2053] = 9'd57;    
		mem[  2054] = 9'd24;    
		mem[  2055] = 9'd46;    
		mem[  2056] = 9'd24;    
		mem[  2057] = 9'd21;    
		mem[  2058] = 9'd21;    
		mem[  2059] = 9'd46;    
		mem[  2060] = 9'd15;    
		mem[  2061] = 9'd32;    
		mem[  2062] = 9'd49;    
		mem[  2063] = 9'd46;    
		mem[  2064] = 9'd24;    
		mem[  2065] = 9'd23;    
		mem[  2066] = 9'd44;    
		mem[  2067] = 9'd46;    
		mem[  2068] = 9'd49;    
		mem[  2069] = 9'd9;    
		mem[  2070] = 9'd10;    
		mem[  2071] = 9'd24;    
		mem[  2072] = 9'd49;    
		mem[  2073] = 9'd43;    
		mem[  2074] = 9'd49;    
		mem[  2075] = 9'd26;    
		mem[  2076] = 9'd9;    
		mem[  2077] = 9'd8;    
		mem[  2078] = 9'd50;    
		mem[  2079] = 9'd21;    
		mem[  2080] = 9'd69;    
		mem[  2081] = 9'd23;    
		mem[  2082] = 9'd71;    
		mem[  2083] = 9'd443;    
		mem[  2084] = 9'd21;    
		mem[  2085] = 9'd80;    
		mem[  2086] = 9'd60;    
		mem[  2087] = 9'd20;    
		mem[  2088] = 9'd80;    
		mem[  2089] = 9'd67;    
		mem[  2090] = 9'd95;    
		mem[  2091] = 9'd48;    
		mem[  2092] = 9'd20;    
		mem[  2093] = 9'd24;    
		mem[  2094] = 9'd49;    
		mem[  2095] = 9'd23;    
		mem[  2096] = 9'd67;    
		mem[  2097] = 9'd22;    
		mem[  2098] = 9'd23;    
		mem[  2099] = 9'd49;    
		mem[  2100] = 9'd47;    
		mem[  2101] = 9'd21;    
		mem[  2102] = 9'd23;    
		mem[  2103] = 9'd48;    
		mem[  2104] = 9'd24;    
		mem[  2105] = 9'd11;    
		mem[  2106] = 9'd56;    
		mem[  2107] = 9'd23;    
		mem[  2108] = 9'd70;    
		mem[  2109] = 9'd42;    
		mem[  2110] = 9'd24;    
		mem[  2111] = 9'd10;    
		mem[  2112] = 9'd10;    
		mem[  2113] = 9'd43;    
		mem[  2114] = 9'd44;    
		mem[  2115] = 9'd45;    
		mem[  2116] = 9'd20;    
		mem[  2117] = 9'd22;    
		mem[  2118] = 9'd44;    
		mem[  2119] = 9'd42;    
		mem[  2120] = 9'd44;    
		mem[  2121] = 9'd21;    
		mem[  2122] = 9'd22;    
		mem[  2123] = 9'd22;    
		mem[  2124] = 9'd22;    
		mem[  2125] = 9'd22;    
		mem[  2126] = 9'd22;    
		mem[  2127] = 9'd22;    
		mem[  2128] = 9'd22;    
		mem[  2129] = 9'd22;    
		mem[  2130] = 9'd21;    
		mem[  2131] = 9'd23;    
		mem[  2132] = 9'd21;    
		mem[  2133] = 9'd22;    
		mem[  2134] = 9'd22;    
		mem[  2135] = 9'd54;    
		mem[  2136] = 9'd31;    
		mem[  2137] = 9'd45;    
		mem[  2138] = 9'd44;    
		mem[  2139] = 9'd21;    
		mem[  2140] = 9'd21;    
		mem[  2141] = 9'd43;    
		mem[  2142] = 9'd43;    
		mem[  2143] = 9'd11;    
		mem[  2144] = 9'd36;    
		mem[  2145] = 9'd23;    
		mem[  2146] = 9'd52;    
		mem[  2147] = 9'd12;    
		mem[  2148] = 9'd44;    
		mem[  2149] = 9'd20;    
		mem[  2150] = 9'd22;    
		mem[  2151] = 9'd22;    
		mem[  2152] = 9'd21;    
		mem[  2153] = 9'd46;    
		mem[  2154] = 9'd44;    
		mem[  2155] = 9'd32;    
		mem[  2156] = 9'd53;    
		mem[  2157] = 9'd45;    
		mem[  2158] = 9'd20;    
		mem[  2159] = 9'd65;    
		mem[  2160] = 9'd44;    
		mem[  2161] = 9'd11;    
		mem[  2162] = 9'd33;    
		mem[  2163] = 9'd34;    
		mem[  2164] = 9'd45;    
		mem[  2165] = 9'd10;    
		mem[  2166] = 9'd43;    
		mem[  2167] = 9'd21;    
		mem[  2168] = 9'd20;    
		mem[  2169] = 9'd24;    
		mem[  2170] = 9'd20;    
		mem[  2171] = 9'd46;    
		mem[  2172] = 9'd43;    
		mem[  2173] = 9'd18;    
		mem[  2174] = 9'd23;    
		mem[  2175] = 9'd46;    
		mem[  2176] = 9'd44;    
		mem[  2177] = 9'd21;    
		mem[  2178] = 9'd64;    
		mem[  2179] = 9'd23;    
		mem[  2180] = 9'd21;    
		mem[  2181] = 9'd20;    
		mem[  2182] = 9'd23;    
		mem[  2183] = 9'd43;    
		mem[  2184] = 9'd44;    
		mem[  2185] = 9'd45;    
		mem[  2186] = 9'd22;    
		mem[  2187] = 9'd20;    
		mem[  2188] = 9'd25;    
		mem[  2189] = 9'd20;    
		mem[  2190] = 9'd45;    
		mem[  2191] = 9'd19;    
		mem[  2192] = 9'd23;    
		mem[  2193] = 9'd21;    
		mem[  2194] = 9'd21;    
		mem[  2195] = 9'd23;    
		mem[  2196] = 9'd23;    
		mem[  2197] = 9'd44;    
		mem[  2198] = 9'd23;    
		mem[  2199] = 9'd9;    
		mem[  2200] = 9'd8;    
		mem[  2201] = 9'd45;    
		mem[  2202] = 9'd45;    
		mem[  2203] = 9'd20;    
		mem[  2204] = 9'd22;    
		mem[  2205] = 9'd43;    
		mem[  2206] = 9'd43;    
		mem[  2207] = 9'd46;    
		mem[  2208] = 9'd23;    
		mem[  2209] = 9'd10;    
		mem[  2210] = 9'd8;    
		mem[  2211] = 9'd35;    
		mem[  2212] = 9'd11;    
		mem[  2213] = 9'd44;    
		mem[  2214] = 9'd20;    
		mem[  2215] = 9'd22;    
		mem[  2216] = 9'd23;    
		mem[  2217] = 9'd20;    
		mem[  2218] = 9'd45;    
		mem[  2219] = 9'd44;    
		mem[  2220] = 9'd42;    
		mem[  2221] = 9'd24;    
		mem[  2222] = 9'd21;    
		mem[  2223] = 9'd44;    
		mem[  2224] = 9'd21;    
		mem[  2225] = 9'd21;    
		mem[  2226] = 9'd43;    
		mem[  2227] = 9'd25;    
		mem[  2228] = 9'd19;    
		mem[  2229] = 9'd21;    
		mem[  2230] = 9'd23;    
		mem[  2231] = 9'd35;    
		mem[  2232] = 9'd44;    
		mem[  2233] = 9'd10;    
		mem[  2234] = 9'd43;    
		mem[  2235] = 9'd21;    
		mem[  2236] = 9'd20;    
		mem[  2237] = 9'd25;    
		mem[  2238] = 9'd19;    
		mem[  2239] = 9'd47;    
		mem[  2240] = 9'd43;    
		mem[  2241] = 9'd17;    
		mem[  2242] = 9'd23;    
		mem[  2243] = 9'd46;    
		mem[  2244] = 9'd44;    
		mem[  2245] = 9'd22;    
		mem[  2246] = 9'd63;    
		mem[  2247] = 9'd44;    
		mem[  2248] = 9'd20;    
		mem[  2249] = 9'd23;    
		mem[  2250] = 9'd42;    
		mem[  2251] = 9'd45;    
		mem[  2252] = 9'd46;    
		mem[  2253] = 9'd27;    
		mem[  2254] = 9'd11;    
		mem[  2255] = 9'd59;    
		mem[  2256] = 9'd23;    
		mem[  2257] = 9'd75;    
		mem[  2258] = 9'd51;    
		mem[  2259] = 9'd45;    
		mem[  2260] = 9'd53;    
		mem[  2261] = 9'd21;    
		mem[  2262] = 9'd25;    
		mem[  2263] = 9'd37;    
		mem[  2264] = 9'd14;    
		mem[  2265] = 9'd48;    
		mem[  2266] = 9'd46;    
		mem[  2267] = 9'd51;    
		mem[  2268] = 9'd24;    
		mem[  2269] = 9'd75;    
		mem[  2270] = 9'd49;    
		mem[  2271] = 9'd20;    
		mem[  2272] = 9'd24;    
		mem[  2273] = 9'd49;    
		mem[  2274] = 9'd23;    
		mem[  2275] = 9'd67;    
		mem[  2276] = 9'd22;    
		mem[  2277] = 9'd23;    
		mem[  2278] = 9'd49;    
		mem[  2279] = 9'd47;    
		mem[  2280] = 9'd21;    
		mem[  2281] = 9'd23;    
		mem[  2282] = 9'd48;    
		mem[  2283] = 9'd24;    
		mem[  2284] = 9'd11;    
		mem[  2285] = 9'd8;    
		mem[  2286] = 9'd48;    
		mem[  2287] = 9'd23;    
		mem[  2288] = 9'd71;    
		mem[  2289] = 9'd46;    
		mem[  2290] = 9'd23;    
		mem[  2291] = 9'd22;    
		mem[  2292] = 9'd45;    
		mem[  2293] = 9'd47;    
		mem[  2294] = 9'd23;    
		mem[  2295] = 9'd23;    
		mem[  2296] = 9'd23;    
		mem[  2297] = 9'd24;    
		mem[  2298] = 9'd23;    
		mem[  2299] = 9'd23;    
		mem[  2300] = 9'd24;    
		mem[  2301] = 9'd22;    
		mem[  2302] = 9'd24;    
		mem[  2303] = 9'd23;    
		mem[  2304] = 9'd23;    
		mem[  2305] = 9'd23;    
		mem[  2306] = 9'd24;    
		mem[  2307] = 9'd67;    
		mem[  2308] = 9'd49;    
		mem[  2309] = 9'd35;    
		mem[  2310] = 9'd8;    
		mem[  2311] = 9'd51;    
		mem[  2312] = 9'd20;    
		mem[  2313] = 9'd69;    
		mem[  2314] = 9'd22;    
		mem[  2315] = 9'd72;    
		mem[  2316] = 9'd45;    
		mem[  2317] = 9'd26;    
		mem[  2318] = 9'd9;    
		mem[  2319] = 9'd12;    
		mem[  2320] = 9'd45;    
		mem[  2321] = 9'd47;    
		mem[  2322] = 9'd48;    
		mem[  2323] = 9'd21;    
		mem[  2324] = 9'd23;    
		mem[  2325] = 9'd47;    
		mem[  2326] = 9'd44;    
		mem[  2327] = 9'd49;    
		mem[  2328] = 9'd44;    
		mem[  2329] = 9'd49;    
		mem[  2330] = 9'd23;    
		mem[  2331] = 9'd68;    
		mem[  2332] = 9'd23;    
		mem[  2333] = 9'd71;    
		mem[  2334] = 9'd19;    
		mem[  2335] = 9'd25;    
		mem[  2336] = 9'd47;    
		mem[  2337] = 9'd45;    
		mem[  2338] = 9'd48;    
		mem[  2339] = 9'd47;    
		mem[  2340] = 9'd22;    
		mem[  2341] = 9'd23;    
		mem[  2342] = 9'd46;    
		mem[  2343] = 9'd46;    
		mem[  2344] = 9'd23;    
		mem[  2345] = 9'd23;    
		mem[  2346] = 9'd24;    
		mem[  2347] = 9'd23;    
		mem[  2348] = 9'd23;    
		mem[  2349] = 9'd23;    
		mem[  2350] = 9'd23;    
		mem[  2351] = 9'd23;    
		mem[  2352] = 9'd23;    
		mem[  2353] = 9'd23;    
		mem[  2354] = 9'd24;    
		mem[  2355] = 9'd23;    
		mem[  2356] = 9'd23;    
		mem[  2357] = 9'd23;    
		mem[  2358] = 9'd23;    
		mem[  2359] = 9'd22;    
		mem[  2360] = 9'd58;    
		mem[  2361] = 9'd27;    
		mem[  2362] = 9'd82;    
		mem[  2363] = 9'd56;    
		mem[  2364] = 9'd24;    
		mem[  2365] = 9'd27;    
		mem[  2366] = 9'd59;    
		mem[  2367] = 9'd25;    
		mem[  2368] = 9'd78;    
		mem[  2369] = 9'd15;    
		mem[  2370] = 9'd42;    
		mem[  2371] = 9'd55;    
		mem[  2372] = 9'd57;    
		mem[  2373] = 9'd31;    
		mem[  2374] = 9'd10;    
		mem[  2375] = 9'd40;    
		mem[  2376] = 9'd28;    
		mem[  2377] = 9'd51;    
		mem[  2378] = 9'd29;    
		mem[  2379] = 9'd10;    
		mem[  2380] = 9'd14;    
		mem[  2381] = 9'd50;    
		mem[  2382] = 9'd51;    
		mem[  2383] = 9'd54;    
		mem[  2384] = 9'd48;    
		mem[  2385] = 9'd56;    
		mem[  2386] = 9'd10;    
		mem[  2387] = 9'd13;    
		mem[  2388] = 9'd24;    
		mem[  2389] = 9'd51;    
		mem[  2390] = 9'd15;    
		mem[  2391] = 9'd38;    
		mem[  2392] = 9'd53;    
		mem[  2393] = 9'd53;    
		mem[  2394] = 9'd13;    
		mem[  2395] = 9'd10;    
		mem[  2396] = 9'd26;    
		mem[  2397] = 9'd54;    
		mem[  2398] = 9'd52;    
		mem[  2399] = 9'd51;    
		mem[  2400] = 9'd26;    
		mem[  2401] = 9'd25;    
		mem[  2402] = 9'd26;    
		mem[  2403] = 9'd25;    
		mem[  2404] = 9'd26;    
		mem[  2405] = 9'd25;    
		mem[  2406] = 9'd26;    
		mem[  2407] = 9'd26;    
		mem[  2408] = 9'd26;    
		mem[  2409] = 9'd25;    
		mem[  2410] = 9'd105;    
		mem[  2411] = 9'd48;    
		mem[  2412] = 9'd56;    
		mem[  2413] = 9'd48;    
		mem[  2414] = 9'd56;    
		mem[  2415] = 9'd48;    
		mem[  2416] = 9'd55;    
		mem[  2417] = 9'd48;    
		mem[  2418] = 9'd55;    
		mem[  2419] = 9'd48;    
		mem[  2420] = 9'd55;    
		mem[  2421] = 9'd48;    
		mem[  2422] = 9'd55;    
		mem[  2423] = 9'd49;    
		mem[  2424] = 9'd55;    
		mem[  2425] = 9'd48;    
		mem[  2426] = 9'd55;    
		mem[  2427] = 9'd48;    
		mem[  2428] = 9'd55;    
		mem[  2429] = 9'd48;    
		mem[  2430] = 9'd55;    
		mem[  2431] = 9'd49;    
		mem[  2432] = 9'd54;    
		mem[  2433] = 9'd49;    
		mem[  2434] = 9'd54;    
		mem[  2435] = 9'd49;    
		mem[  2436] = 9'd55;    
		mem[  2437] = 9'd51;    
		mem[  2438] = 9'd27;    
		mem[  2439] = 9'd24;    
		mem[  2440] = 9'd26;    
		mem[  2441] = 9'd25;    
		mem[  2442] = 9'd26;    
		mem[  2443] = 9'd26;    
		mem[  2444] = 9'd25;    
		mem[  2445] = 9'd26;    
		mem[  2446] = 9'd26;    
		mem[  2447] = 9'd26;    
		mem[  2448] = 9'd25;    
		mem[  2449] = 9'd26;    
		mem[  2450] = 9'd26;    
		mem[  2451] = 9'd92;    
		mem[  2452] = 9'd58;    
		mem[  2453] = 9'd64;    
		mem[  2454] = 9'd58;    
		mem[  2455] = 9'd66;    
		mem[  2456] = 9'd57;    
		mem[  2457] = 9'd65;    
		mem[  2458] = 9'd58;    
		mem[  2459] = 9'd65;    
		mem[  2460] = 9'd58;    
		mem[  2461] = 9'd64;    
		mem[  2462] = 9'd58;    
		mem[  2463] = 9'd65;    
		mem[  2464] = 9'd58;    
		mem[  2465] = 9'd64;    
		mem[  2466] = 9'd58;    
		mem[  2467] = 9'd65;    
		mem[  2468] = 9'd58;    
		mem[  2469] = 9'd64;    
		mem[  2470] = 9'd58;    
		mem[  2471] = 9'd65;    
		mem[  2472] = 9'd58;    
		mem[  2473] = 9'd64;    
		mem[  2474] = 9'd61;    
		mem[  2475] = 9'd32;    
		mem[  2476] = 9'd28;    
		mem[  2477] = 9'd32;    
		mem[  2478] = 9'd29;    
		mem[  2479] = 9'd31;    
		mem[  2480] = 9'd30;    
		mem[  2481] = 9'd31;    
		mem[  2482] = 9'd30;    
		mem[  2483] = 9'd31;    
		mem[  2484] = 9'd31;    
		mem[  2485] = 9'd30;    
		mem[  2486] = 9'd94;    
		mem[  2487] = 9'd59;    
		mem[  2488] = 9'd63;    
		mem[  2489] = 9'd60;    
		mem[  2490] = 9'd64;    
		mem[  2491] = 9'd32;    
		mem[  2492] = 9'd10;    
		mem[  2493] = 9'd19;    
		mem[  2494] = 9'd58;    
		mem[  2495] = 9'd64;    
		mem[  2496] = 9'd59;    
		mem[  2497] = 9'd60;    
		mem[  2498] = 9'd32;    
		mem[  2499] = 9'd64;    
		mem[  2500] = 9'd31;    
		mem[  2501] = 9'd13;    
		mem[  2502] = 9'd15;    
		mem[  2503] = 9'd93;    
		mem[  2504] = 9'd36;    
		mem[  2505] = 9'd11;    
		mem[  2506] = 9'd11;    
		mem[  2507] = 9'd66;    
		mem[  2508] = 9'd33;    
		mem[  2509] = 9'd24;    
		mem[  2510] = 9'd65;    
		mem[  2511] = 9'd25;    
		mem[  2512] = 9'd34;    
		mem[  2513] = 9'd62;    
		mem[  2514] = 9'd61;    
		mem[  2515] = 9'd63;    
		mem[  2516] = 9'd31;    
		mem[  2517] = 9'd30;    
		mem[  2518] = 9'd29;    
		mem[  2519] = 9'd31;    
		mem[  2520] = 9'd31;    
		mem[  2521] = 9'd30;    
		mem[  2522] = 9'd31;    
		mem[  2523] = 9'd30;    
		mem[  2524] = 9'd31;    
		mem[  2525] = 9'd30;    
		mem[  2526] = 9'd32;    
		mem[  2527] = 9'd30;    
		mem[  2528] = 9'd31;    
		mem[  2529] = 9'd30;    
		mem[  2530] = 9'd54;    
		mem[  2531] = 9'd59;    
		mem[  2532] = 9'd26;    
		mem[  2533] = 9'd12;    
		mem[  2534] = 9'd71;    
		mem[  2535] = 9'd13;    
		mem[  2536] = 9'd11;    
		mem[  2537] = 9'd30;    
		mem[  2538] = 9'd51;    
		mem[  2539] = 9'd59;    
		mem[  2540] = 9'd26;    
		mem[  2541] = 9'd14;    
		mem[  2542] = 9'd9;    
		mem[  2543] = 9'd60;    
		mem[  2544] = 9'd26;    
		mem[  2545] = 9'd28;    
		mem[  2546] = 9'd82;    
		mem[  2547] = 9'd28;    
		mem[  2548] = 9'd26;    
		mem[  2549] = 9'd24;    
		mem[  2550] = 9'd57;    
		mem[  2551] = 9'd26;    
		mem[  2552] = 9'd13;    
		mem[  2553] = 9'd26;    
		mem[  2554] = 9'd9;    
		mem[  2555] = 9'd25;    
		mem[  2556] = 9'd56;    
		mem[  2557] = 9'd49;    
		mem[  2558] = 9'd52;    
		mem[  2559] = 9'd52;    
		mem[  2560] = 9'd50;    
		mem[  2561] = 9'd53;    
		mem[  2562] = 9'd53;    
		mem[  2563] = 9'd24;    
		mem[  2564] = 9'd79;    
		mem[  2565] = 9'd24;    
		mem[  2566] = 9'd27;    
		mem[  2567] = 9'd50;    
		mem[  2568] = 9'd54;    
		mem[  2569] = 9'd26;    
		mem[  2570] = 9'd23;    
		mem[  2571] = 9'd54;    
		mem[  2572] = 9'd27;    
		mem[  2573] = 9'd21;    
		mem[  2574] = 9'd28;    
		mem[  2575] = 9'd24;    
		mem[  2576] = 9'd55;    
		mem[  2577] = 9'd51;    
		mem[  2578] = 9'd50;    
		mem[  2579] = 9'd53;    
		mem[  2580] = 9'd25;    
		mem[  2581] = 9'd25;    
		mem[  2582] = 9'd52;    
		mem[  2583] = 9'd54;    
		mem[  2584] = 9'd24;    
		mem[  2585] = 9'd24;    
		mem[  2586] = 9'd29;    
		mem[  2587] = 9'd26;    
		mem[  2588] = 9'd24;    
		mem[  2589] = 9'd27;    
		mem[  2590] = 9'd50;    
		mem[  2591] = 9'd28;    
		mem[  2592] = 9'd26;    
		mem[  2593] = 9'd27;    
		mem[  2594] = 9'd22;    
		mem[  2595] = 9'd54;    
		mem[  2596] = 9'd28;    
		mem[  2597] = 9'd21;    
		mem[  2598] = 9'd27;    
		mem[  2599] = 9'd15;    
		mem[  2600] = 9'd10;    
		mem[  2601] = 9'd53;    
		mem[  2602] = 9'd52;    
		mem[  2603] = 9'd50;    
		mem[  2604] = 9'd30;    
		mem[  2605] = 9'd23;    
		mem[  2606] = 9'd51;    
		mem[  2607] = 9'd51;    
		mem[  2608] = 9'd29;    
		mem[  2609] = 9'd24;    
		mem[  2610] = 9'd25;    
		mem[  2611] = 9'd25;    
		mem[  2612] = 9'd25;    
		mem[  2613] = 9'd27;    
		mem[  2614] = 9'd26;    
		mem[  2615] = 9'd26;    
		mem[  2616] = 9'd26;    
		mem[  2617] = 9'd26;    
		mem[  2618] = 9'd26;    
		mem[  2619] = 9'd25;    
		mem[  2620] = 9'd26;    
		mem[  2621] = 9'd26;    
		mem[  2622] = 9'd26;    
		mem[  2623] = 9'd26;    
		mem[  2624] = 9'd26;    
		mem[  2625] = 9'd25;    
		mem[  2626] = 9'd27;    
		mem[  2627] = 9'd25;    
		mem[  2628] = 9'd26;    
		mem[  2629] = 9'd25;    
		mem[  2630] = 9'd27;    
		mem[  2631] = 9'd25;    
		mem[  2632] = 9'd26;    
		mem[  2633] = 9'd26;    
		mem[  2634] = 9'd26;    
		mem[  2635] = 9'd25;    
		mem[  2636] = 9'd26;    
		mem[  2637] = 9'd26;    
		mem[  2638] = 9'd26;    
		mem[  2639] = 9'd25;    
		mem[  2640] = 9'd27;    
		mem[  2641] = 9'd52;    
		mem[  2642] = 9'd27;    
		mem[  2643] = 9'd48;    
		mem[  2644] = 9'd56;    
		mem[  2645] = 9'd24;    
		mem[  2646] = 9'd15;    
		mem[  2647] = 9'd7;    
		mem[  2648] = 9'd56;    
		mem[  2649] = 9'd25;    
		mem[  2650] = 9'd25;    
		mem[  2651] = 9'd78;    
		mem[  2652] = 9'd27;    
		mem[  2653] = 9'd26;    
		mem[  2654] = 9'd22;    
		mem[  2655] = 9'd55;    
		mem[  2656] = 9'd26;    
		mem[  2657] = 9'd10;    
		mem[  2658] = 9'd14;    
		mem[  2659] = 9'd79;    
		mem[  2660] = 9'd26;    
		mem[  2661] = 9'd27;    
		mem[  2662] = 9'd21;    
		mem[  2663] = 9'd55;    
		mem[  2664] = 9'd26;    
		mem[  2665] = 9'd12;    
		mem[  2666] = 9'd12;    
		mem[  2667] = 9'd12;    
		mem[  2668] = 9'd66;    
		mem[  2669] = 9'd27;    
		mem[  2670] = 9'd28;    
		mem[  2671] = 9'd20;    
		mem[  2672] = 9'd55;    
		mem[  2673] = 9'd27;    
		mem[  2674] = 9'd13;    
		mem[  2675] = 9'd34;    
		mem[  2676] = 9'd25;    
		mem[  2677] = 9'd28;    
		mem[  2678] = 9'd28;    
		mem[  2679] = 9'd49;    
		mem[  2680] = 9'd54;    
		mem[  2681] = 9'd27;    
		mem[  2682] = 9'd15;    
		mem[  2683] = 9'd23;    
		mem[  2684] = 9'd10;    
		mem[  2685] = 9'd25;    
		mem[  2686] = 9'd34;    
		mem[  2687] = 9'd33;    
		mem[  2688] = 9'd30;    
		mem[  2689] = 9'd30;    
		mem[  2690] = 9'd67;    
		mem[  2691] = 9'd34;    
		mem[  2692] = 9'd29;    
		mem[  2693] = 9'd36;    
		mem[  2694] = 9'd34;    
		mem[  2695] = 9'd30;    
		mem[  2696] = 9'd30;    
		mem[  2697] = 9'd67;    
		mem[  2698] = 9'd33;    
		mem[  2699] = 9'd30;    
		mem[  2700] = 9'd36;    
		mem[  2701] = 9'd33;    
		mem[  2702] = 9'd31;    
		mem[  2703] = 9'd30;    
		mem[  2704] = 9'd67;    
		mem[  2705] = 9'd33;    
		mem[  2706] = 9'd16;    
		mem[  2707] = 9'd12;    
		mem[  2708] = 9'd32;    
		mem[  2709] = 9'd33;    
		mem[  2710] = 9'd30;    
		mem[  2711] = 9'd17;    
		mem[  2712] = 9'd11;    
		mem[  2713] = 9'd34;    
		mem[  2714] = 9'd30;    
		mem[  2715] = 9'd59;    
		mem[  2716] = 9'd63;    
		mem[  2717] = 9'd32;    
		mem[  2718] = 9'd28;    
		mem[  2719] = 9'd63;    
		mem[  2720] = 9'd30;    
		mem[  2721] = 9'd30;    
		mem[  2722] = 9'd61;    
		mem[  2723] = 9'd62;    
		mem[  2724] = 9'd61;    
		mem[  2725] = 9'd62;    
		mem[  2726] = 9'd33;    
		mem[  2727] = 9'd28;    
		mem[  2728] = 9'd31;    
		mem[  2729] = 9'd30;    
		mem[  2730] = 9'd31;    
		mem[  2731] = 9'd30;    
		mem[  2732] = 9'd30;    
		mem[  2733] = 9'd31;    
		mem[  2734] = 9'd30;    
		mem[  2735] = 9'd31;    
		mem[  2736] = 9'd30;    
		mem[  2737] = 9'd31;    
		mem[  2738] = 9'd31;    
		mem[  2739] = 9'd30;    
		mem[  2740] = 9'd31;    
		mem[  2741] = 9'd31;    
		mem[  2742] = 9'd31;    
		mem[  2743] = 9'd30;    
		mem[  2744] = 9'd31;    
		mem[  2745] = 9'd30;    
		mem[  2746] = 9'd31;    
		mem[  2747] = 9'd31;    
		mem[  2748] = 9'd29;    
		mem[  2749] = 9'd33;    
		mem[  2750] = 9'd59;    
		mem[  2751] = 9'd63;    
		mem[  2752] = 9'd63;    
		mem[  2753] = 9'd31;    
		mem[  2754] = 9'd30;    
		mem[  2755] = 9'd59;    
		mem[  2756] = 9'd63;    
		mem[  2757] = 9'd62;    
		mem[  2758] = 9'd31;    
		mem[  2759] = 9'd30;    
		mem[  2760] = 9'd59;    
		mem[  2761] = 9'd62;    
		mem[  2762] = 9'd63;    
		mem[  2763] = 9'd31;    
		mem[  2764] = 9'd30;    
		mem[  2765] = 9'd59;    
		mem[  2766] = 9'd63;    
		mem[  2767] = 9'd62;    
		mem[  2768] = 9'd31;    
		mem[  2769] = 9'd30;    
		mem[  2770] = 9'd59;    
		mem[  2771] = 9'd63;    
		mem[  2772] = 9'd62;    
		mem[  2773] = 9'd31;    
		mem[  2774] = 9'd30;    
		mem[  2775] = 9'd60;    
		mem[  2776] = 9'd62;    
		mem[  2777] = 9'd62;    
		mem[  2778] = 9'd31;    
		mem[  2779] = 9'd30;    
		mem[  2780] = 9'd60;    
		mem[  2781] = 9'd62;    
		mem[  2782] = 9'd62;    
		mem[  2783] = 9'd31;    
		mem[  2784] = 9'd30;    
		mem[  2785] = 9'd60;    
		mem[  2786] = 9'd62;    
		mem[  2787] = 9'd62;    
		mem[  2788] = 9'd31;    
		mem[  2789] = 9'd30;    
		mem[  2790] = 9'd60;    
		mem[  2791] = 9'd62;    
		mem[  2792] = 9'd62;    
		mem[  2793] = 9'd31;    
		mem[  2794] = 9'd30;    
		mem[  2795] = 9'd60;    
		mem[  2796] = 9'd62;    
		mem[  2797] = 9'd62;    
		mem[  2798] = 9'd31;    
		mem[  2799] = 9'd30;    
		mem[  2800] = 9'd60;    
		mem[  2801] = 9'd62;    
		mem[  2802] = 9'd62;    
		mem[  2803] = 9'd31;    
		mem[  2804] = 9'd30;    
		mem[  2805] = 9'd60;    
		mem[  2806] = 9'd62;    
		mem[  2807] = 9'd63;    
		mem[  2808] = 9'd31;    
		mem[  2809] = 9'd30;    
		mem[  2810] = 9'd59;    
		mem[  2811] = 9'd62;    
		mem[  2812] = 9'd63;    
		mem[  2813] = 9'd31;    
		mem[  2814] = 9'd30;    
		mem[  2815] = 9'd59;    
		mem[  2816] = 9'd62;    
		mem[  2817] = 9'd63;    
		mem[  2818] = 9'd31;    
		mem[  2819] = 9'd30;    
		mem[  2820] = 9'd59;    
		mem[  2821] = 9'd62;    
		mem[  2822] = 9'd62;    
		mem[  2823] = 9'd32;    
		mem[  2824] = 9'd30;    
		mem[  2825] = 9'd59;    
		mem[  2826] = 9'd62;    
		mem[  2827] = 9'd63;    
		mem[  2828] = 9'd31;    
		mem[  2829] = 9'd30;    
		mem[  2830] = 9'd59;    
		mem[  2831] = 9'd62;    
		mem[  2832] = 9'd63;    
		mem[  2833] = 9'd31;    
		mem[  2834] = 9'd30;    
		mem[  2835] = 9'd59;    
		mem[  2836] = 9'd62;    
		mem[  2837] = 9'd511;    
		mem[  2838] = 9'd511;    
	end
	
endmodule

